-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 21 2024 23:56:49

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    masterreset : in std_logic;
    led4 : out std_logic;
    lcol3 : out std_logic;
    led5 : out std_logic;
    lcol2 : out std_logic;
    led6 : out std_logic;
    led2 : out std_logic;
    lcol1 : out std_logic;
    deldn : in std_logic;
    cpuclk : out std_logic;
    apureset : out std_logic;
    altreset : in std_logic;
    led7 : out std_logic;
    led3 : out std_logic;
    lcol4 : out std_logic;
    delup : in std_logic;
    cpureset : out std_logic;
    apusync : in std_logic;
    PACKAGEPIN : in std_logic;
    led8 : out std_logic;
    led1 : out std_logic;
    consolereset : in std_logic;
    apuclk : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2196\ : std_logic;
signal \arse.un1_io_0_1_g\ : std_logic;
signal \top_pll_nrtthrth.PLLOUTCORE\ : std_logic;
signal \GNDG0\ : std_logic;
signal \arse.divseven.io_0_D_IN_0\ : std_logic;
signal \VCCG0\ : std_logic;
signal masterreset_c_i : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \debounceup.un3_counter_1_cry_1\ : std_logic;
signal \debounceup.un3_counter_1_cry_2\ : std_logic;
signal \debounceup.un3_counter_1_cry_3\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \arses.un2_counter_cry_1\ : std_logic;
signal \arses.un2_counter_cry_2\ : std_logic;
signal \arses.un2_counter_cry_3\ : std_logic;
signal \arses.un2_counter_cry_4\ : std_logic;
signal \arses.un2_counter_cry_5\ : std_logic;
signal \arses.un2_counter_cry_6\ : std_logic;
signal \arses.un2_counter_cry_7\ : std_logic;
signal \arses.un2_counter_cry_8\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \arses.un2_counter_cry_9\ : std_logic;
signal \arses.un2_counter_cry_10\ : std_logic;
signal \arses.un2_counter_cry_11\ : std_logic;
signal \arses.un2_counter_cry_12\ : std_logic;
signal \arses.un2_counter_cry_13\ : std_logic;
signal lcol4_c : std_logic;
signal \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\ : std_logic;
signal \debounceup.counterZ0Z_3\ : std_logic;
signal \debounceup.counter19_2_cascade_\ : std_logic;
signal \debounceup.counter_RNO_0_0_2\ : std_logic;
signal \debounceup.counter19_cascade_\ : std_logic;
signal \debounceup.counterZ0Z_2\ : std_logic;
signal \debounceup.counterZ0Z_4\ : std_logic;
signal \debounceup.counter19_2\ : std_logic;
signal \dig2.m18_bm_cascade_\ : std_logic;
signal leds_1_i_1 : std_logic;
signal \arses.counterZ0Z_7\ : std_logic;
signal \arses.counterZ0Z_6\ : std_logic;
signal \arses.counterZ0Z_5\ : std_logic;
signal \arses.counterZ0Z_8\ : std_logic;
signal \arses.counterZ0Z_3\ : std_logic;
signal \arses.counterZ0Z_2\ : std_logic;
signal \arses.counterZ0Z_4\ : std_logic;
signal \arses.un1_counterlto4_2_cascade_\ : std_logic;
signal \arses.un1_counterlto8_2\ : std_logic;
signal \arses.counterZ0Z_11\ : std_logic;
signal \arses.counterZ0Z_10\ : std_logic;
signal \arses.un1_counterlt11_cascade_\ : std_logic;
signal \arses.counterZ0Z_9\ : std_logic;
signal \arses.counterZ0Z_14\ : std_logic;
signal \arses.counterZ0Z_13\ : std_logic;
signal \arses.un1_counterlt13_0_cascade_\ : std_logic;
signal \arses.counterZ0Z_12\ : std_logic;
signal \arses_counter8_cascade_\ : std_logic;
signal \arses.clock_out_RNIR6ERZ0Z_0\ : std_logic;
signal \arses.counterZ0Z_1\ : std_logic;
signal \arses.counterZ0Z_0\ : std_logic;
signal lcol3_c : std_logic;
signal \dig2.m13_am_cascade_\ : std_logic;
signal \dig2.leds_17_i_0_ns_1_1\ : std_logic;
signal \dig2.m18_am\ : std_logic;
signal leds_1_i_3 : std_logic;
signal \dig2.m13_bm\ : std_logic;
signal \dig2.N_42\ : std_logic;
signal \dig2.m69_am\ : std_logic;
signal \dig2.m69_bm\ : std_logic;
signal leds_1_i_0_2 : std_logic;
signal \dig2.N_78\ : std_logic;
signal \dig2.N_76\ : std_logic;
signal leds_1_i_0_3 : std_logic;
signal \dig2.m39_ns_1_cascade_\ : std_logic;
signal \dig2.N_40\ : std_logic;
signal \dig2.i3_mux\ : std_logic;
signal \dig2.N_59\ : std_logic;
signal \dig2.leds_17_i_ns_1_2\ : std_logic;
signal consolereset_c : std_logic;
signal altreset_c : std_logic;
signal \debounceconsolereset.out_RNOZ0Z_0_cascade_\ : std_logic;
signal \clock_out_RNIR6ER\ : std_logic;
signal \clock_out_RNIR6ER_cascade_\ : std_logic;
signal arses_counter8 : std_logic;
signal slowclk : std_logic;
signal \dig2.m54_am\ : std_logic;
signal leds_1_i_0_1 : std_logic;
signal \dig2.m75_ns_1\ : std_logic;
signal \bfn_20_17_0_\ : std_logic;
signal \debounceconsolereset.counter_RNO_0Z0Z_2\ : std_logic;
signal \debounceconsolereset.un3_counter_1_cry_1\ : std_logic;
signal \debounceconsolereset.un3_counter_1_cry_2\ : std_logic;
signal \debounceconsolereset.un3_counter_1_cry_3\ : std_logic;
signal \debounceconsolereset.counterZ0Z_3\ : std_logic;
signal \debounceconsolereset.counterZ0Z_2\ : std_logic;
signal \debounceconsolereset.counter19_2\ : std_logic;
signal \debounceconsolereset.counterZ0Z_4\ : std_logic;
signal \debounceconsolereset.counterZ0Z_1\ : std_logic;
signal \debounceconsolereset.counter19_2_cascade_\ : std_logic;
signal \debounceconsolereset.counterZ0Z_0\ : std_logic;
signal \debounceconsolereset.counter19\ : std_logic;
signal col_1_1 : std_logic;
signal \dig2.m54_bm\ : std_logic;
signal \dig2.leds_17_i_ns_1_1\ : std_logic;
signal \debounceup.counterZ0Z_0\ : std_logic;
signal \debounceup.counterZ0Z_1\ : std_logic;
signal \dig2.m49_bm\ : std_logic;
signal \dig2.m49_am\ : std_logic;
signal \dig2.m33_am\ : std_logic;
signal \dig2.m33_bm_cascade_\ : std_logic;
signal leds_1_i_2 : std_logic;
signal \dig2.N_25_cascade_\ : std_logic;
signal \dig2.leds_17_i_0_ns_1_2\ : std_logic;
signal \dig2.i2_mux\ : std_logic;
signal lcol1_c : std_logic;
signal \colZ0Z_1\ : std_logic;
signal \colZ0Z_0\ : std_logic;
signal lcol2_c : std_logic;
signal \debouncedn.counter19_2_cascade_\ : std_logic;
signal \debouncedn.counter19_cascade_\ : std_logic;
signal \bfn_24_17_0_\ : std_logic;
signal \debouncedn.counterZ0Z_2\ : std_logic;
signal \debouncedn.counter_RNO_0_1_2\ : std_logic;
signal \debouncedn.un3_counter_1_cry_1\ : std_logic;
signal \debouncedn.counterZ0Z_3\ : std_logic;
signal \debouncedn.un3_counter_1_cry_2\ : std_logic;
signal \debouncedn.counter19_2\ : std_logic;
signal \debouncedn.un3_counter_1_cry_3\ : std_logic;
signal \debouncedn.counterZ0Z_4\ : std_logic;
signal \debouncedn.counterZ0Z_0\ : std_logic;
signal \debouncedn.counterZ0Z_1\ : std_logic;
signal \debouncedn.counter19\ : std_logic;
signal deldn_c : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bfn_27_10_0_\ : std_logic;
signal \un1_delayConstant_cry_0\ : std_logic;
signal \un1_delayConstant_cry_1\ : std_logic;
signal \un1_delayConstant_cry_2\ : std_logic;
signal \delayConstantZ0Z_4\ : std_logic;
signal \un1_delayConstant_cry_3\ : std_logic;
signal \delayConstantZ0Z_5\ : std_logic;
signal \un1_delayConstant_cry_4\ : std_logic;
signal \delayConstantZ0Z_6\ : std_logic;
signal \un1_delayConstant_cry_5\ : std_logic;
signal \un1_delayConstant_cry_6\ : std_logic;
signal \delayConstantZ0Z_7\ : std_logic;
signal masterreset_c_i_g : std_logic;
signal \olddnZ0\ : std_logic;
signal debounceddn : std_logic;
signal \olddn_RNIEENHZ0_cascade_\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_0\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_3\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_1\ : std_logic;
signal masterreset_c : std_logic;
signal \delayConstant17_i_cascade_\ : std_logic;
signal \un1_delayConstant_cry_0_c_RNOZ0\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_4\ : std_logic;
signal \olddn_RNIM5BHZ0Z1\ : std_logic;
signal \olddn_RNIEENHZ0\ : std_logic;
signal \delayConstant17_i\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_2\ : std_logic;
signal \oldupZ0\ : std_logic;
signal \debounceup.counter19\ : std_logic;
signal delup_c : std_logic;
signal \N_111_g\ : std_logic;
signal debouncedup : std_logic;
signal \PACKAGEPIN_0_c_g\ : std_logic;
signal \bfn_29_7_0_\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_0\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_1\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_2\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_3\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_4\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_5\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_6\ : std_logic;
signal \INVarse.cpuresetcount_0C_net\ : std_logic;
signal \arse.cpuresetoutregZ0\ : std_logic;
signal \INVarse.cpuresetoutregC_net\ : std_logic;
signal \arse.m8_2_cascade_\ : std_logic;
signal \arse.cpuresetcountZ0Z_0\ : std_logic;
signal \arse.cpuresetcountZ0Z_5\ : std_logic;
signal \arse.cpuresetcountZ0Z_1\ : std_logic;
signal \arse.cpuresetcountZ0Z_2\ : std_logic;
signal \arse.m12_2_cascade_\ : std_logic;
signal \arse.cpuresetcountZ0Z_4\ : std_logic;
signal \arse.cpuresetoutreg_1_sqmuxa\ : std_logic;
signal \arse.cpuresetcountZ0Z_7\ : std_logic;
signal \arse.cpuresetcountZ0Z_6\ : std_logic;
signal \arse.cpuresetcountZ0Z_3\ : std_logic;
signal \arse.m4_e_2\ : std_logic;
signal \arse.cpuclkreset_1_sqmuxa\ : std_logic;
signal \INVarse.cpuclkresetC_net\ : std_logic;
signal debouncedconsolereset_i : std_logic;
signal \INVarse.diveight.dout_0C_net\ : std_logic;
signal \delayConstantZ0Z_3\ : std_logic;
signal \arse_diveight_N_123_0_cascade_\ : std_logic;
signal \delayConstantZ0Z_2\ : std_logic;
signal \delayConstantZ0Z_1\ : std_logic;
signal arse_cpuclkreset : std_logic;
signal apusync_c : std_logic;
signal \arse.apusynclatchedZ0\ : std_logic;
signal \INVarse.apusynclatchedC_net\ : std_logic;
signal \arse.diveight.doutZ0Z_0\ : std_logic;
signal \arse.diveight.dout_i_0\ : std_logic;
signal \arse.diveight.dout_i_1\ : std_logic;
signal debouncedconsolereset : std_logic;
signal \arse.apuresetoutregZ0\ : std_logic;
signal \INVarse.apuresetoutregC_net\ : std_logic;
signal arse_diveight_counter_1 : std_logic;
signal arse_diveight_counter_0 : std_logic;
signal \delayConstantZ0Z_0\ : std_logic;
signal arse_diveight_counter_2 : std_logic;
signal \arse.diveight.doutZ0Z_1\ : std_logic;
signal \arse.diveight.cpuclkreset_i\ : std_logic;
signal \arse.divseven.counterZ0Z_1\ : std_logic;
signal \arse.divseven.counterZ0Z_0\ : std_logic;
signal \INVarse.divseven.dout_0C_net\ : std_logic;
signal \arse.divseven.doutZ0Z_0\ : std_logic;
signal \arse.divseven.dout_i_0\ : std_logic;
signal \arse.divseven.counterZ0Z_2\ : std_logic;
signal \PLLOUTCORE_g\ : std_logic;
signal \arse.divseven.doutZ0Z_1\ : std_logic;
signal \arse.divseven.dout_i_1\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PACKAGEPIN_wire\ : std_logic;
signal masterreset_wire : std_logic;
signal led3_wire : std_logic;
signal apuclk_wire : std_logic;
signal cpureset_wire : std_logic;
signal lcol3_wire : std_logic;
signal deldn_wire : std_logic;
signal led2_wire : std_logic;
signal delup_wire : std_logic;
signal led6_wire : std_logic;
signal led8_wire : std_logic;
signal altreset_wire : std_logic;
signal led4_wire : std_logic;
signal apureset_wire : std_logic;
signal lcol4_wire : std_logic;
signal cpuclk_wire : std_logic;
signal led5_wire : std_logic;
signal consolereset_wire : std_logic;
signal lcol2_wire : std_logic;
signal led1_wire : std_logic;
signal apusync_wire : std_logic;
signal led7_wire : std_logic;
signal lcol1_wire : std_logic;
signal \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \PACKAGEPIN_wire\ <= PACKAGEPIN;
    masterreset_wire <= masterreset;
    led3 <= led3_wire;
    apuclk <= apuclk_wire;
    cpureset <= cpureset_wire;
    lcol3 <= lcol3_wire;
    deldn_wire <= deldn;
    led2 <= led2_wire;
    delup_wire <= delup;
    led6 <= led6_wire;
    led8 <= led8_wire;
    altreset_wire <= altreset;
    led4 <= led4_wire;
    apureset <= apureset_wire;
    lcol4 <= lcol4_wire;
    cpuclk <= cpuclk_wire;
    led5 <= led5_wire;
    consolereset_wire <= consolereset;
    lcol2 <= lcol2_wire;
    led1 <= led1_wire;
    apusync_wire <= apusync;
    led7 <= led7_wire;
    lcol1 <= lcol1_wire;
    \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_nrtthrth.top_pll_nrtthrth_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "010",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \top_pll_nrtthrth.PLLOUTCORE\,
            REFERENCECLK => \N__2304\,
            RESETB => \N__4878\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PACKAGEPIN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6028\,
            GLOBALBUFFEROUTPUT => \PACKAGEPIN_0_c_g\
        );

    \PACKAGEPIN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6030\,
            DIN => \N__6029\,
            DOUT => \N__6028\,
            PACKAGEPIN => \PACKAGEPIN_wire\
        );

    \PACKAGEPIN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6030\,
            PADOUT => \N__6029\,
            PADIN => \N__6028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \masterreset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6019\,
            DIN => \N__6018\,
            DOUT => \N__6017\,
            PACKAGEPIN => masterreset_wire
        );

    \masterreset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6019\,
            PADOUT => \N__6018\,
            PADIN => \N__6017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => masterreset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6010\,
            DIN => \N__6009\,
            DOUT => \N__6008\,
            PACKAGEPIN => led3_wire
        );

    \led3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6010\,
            PADOUT => \N__6009\,
            PADIN => \N__6008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2820\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.divseven.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6001\,
            DIN => \N__6000\,
            DOUT => \N__5999\,
            PACKAGEPIN => apuclk_wire
        );

    \arse.divseven.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6001\,
            PADOUT => \N__6000\,
            PADIN => \N__5999\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__5697\,
            OUTPUTENABLE => \N__3832\,
            DIN0 => \arse.divseven.io_0_D_IN_0\,
            DOUT0 => \N__5778\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5738\
        );

    \arse.io_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5992\,
            DIN => \N__5991\,
            DOUT => \N__5990\,
            PACKAGEPIN => cpureset_wire
        );

    \arse.io_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5992\,
            PADOUT => \N__5991\,
            PADIN => \N__5990\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4896\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5748\
        );

    \lcol3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5983\,
            DIN => \N__5982\,
            DOUT => \N__5981\,
            PACKAGEPIN => lcol3_wire
        );

    \lcol3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5983\,
            PADOUT => \N__5982\,
            PADIN => \N__5981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2556\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \deldn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5974\,
            DIN => \N__5973\,
            DOUT => \N__5972\,
            PACKAGEPIN => deldn_wire
        );

    \deldn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5974\,
            PADOUT => \N__5973\,
            PADIN => \N__5972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => deldn_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5965\,
            DIN => \N__5964\,
            DOUT => \N__5963\,
            PACKAGEPIN => led2_wire
        );

    \led2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5965\,
            PADOUT => \N__5964\,
            PADIN => \N__5963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2856\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delup_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5956\,
            DIN => \N__5955\,
            DOUT => \N__5954\,
            PACKAGEPIN => delup_wire
        );

    \delup_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5956\,
            PADOUT => \N__5955\,
            PADIN => \N__5954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delup_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led6_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5947\,
            DIN => \N__5946\,
            DOUT => \N__5945\,
            PACKAGEPIN => led6_wire
        );

    \led6_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5947\,
            PADOUT => \N__5946\,
            PADIN => \N__5945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led8_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5938\,
            DIN => \N__5937\,
            DOUT => \N__5936\,
            PACKAGEPIN => led8_wire
        );

    \led8_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5938\,
            PADOUT => \N__5937\,
            PADIN => \N__5936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \altreset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5929\,
            DIN => \N__5928\,
            DOUT => \N__5927\,
            PACKAGEPIN => altreset_wire
        );

    \altreset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5929\,
            PADOUT => \N__5928\,
            PADIN => \N__5927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => altreset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5920\,
            DIN => \N__5919\,
            DOUT => \N__5918\,
            PACKAGEPIN => led4_wire
        );

    \led4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5920\,
            PADOUT => \N__5919\,
            PADIN => \N__5918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2784\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5911\,
            DIN => \N__5910\,
            DOUT => \N__5909\,
            PACKAGEPIN => apureset_wire
        );

    \arse.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5911\,
            PADOUT => \N__5910\,
            PADIN => \N__5909\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5376\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5744\
        );

    \lcol4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5902\,
            DIN => \N__5901\,
            DOUT => \N__5900\,
            PACKAGEPIN => lcol4_wire
        );

    \lcol4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5902\,
            PADOUT => \N__5901\,
            PADIN => \N__5900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2322\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.diveight.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5893\,
            DIN => \N__5892\,
            DOUT => \N__5891\,
            PACKAGEPIN => cpuclk_wire
        );

    \arse.diveight.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5893\,
            PADOUT => \N__5892\,
            PADIN => \N__5891\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__5430\,
            OUTPUTENABLE => \N__3840\,
            DIN0 => OPEN,
            DOUT0 => \N__5436\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5744\
        );

    \led5_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5884\,
            DIN => \N__5883\,
            DOUT => \N__5882\,
            PACKAGEPIN => led5_wire
        );

    \led5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5884\,
            PADOUT => \N__5883\,
            PADIN => \N__5882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3836\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \consolereset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5875\,
            DIN => \N__5874\,
            DOUT => \N__5873\,
            PACKAGEPIN => consolereset_wire
        );

    \consolereset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5875\,
            PADOUT => \N__5874\,
            PADIN => \N__5873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => consolereset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5866\,
            DIN => \N__5865\,
            DOUT => \N__5864\,
            PACKAGEPIN => lcol2_wire
        );

    \lcol2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5866\,
            PADOUT => \N__5865\,
            PADIN => \N__5864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3405\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5857\,
            DIN => \N__5856\,
            DOUT => \N__5855\,
            PACKAGEPIN => led1_wire
        );

    \led1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5857\,
            PADOUT => \N__5856\,
            PADIN => \N__5855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3819\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \apusync_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5848\,
            DIN => \N__5847\,
            DOUT => \N__5846\,
            PACKAGEPIN => apusync_wire
        );

    \apusync_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5848\,
            PADOUT => \N__5847\,
            PADIN => \N__5846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => apusync_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5839\,
            DIN => \N__5838\,
            DOUT => \N__5837\,
            PACKAGEPIN => led7_wire
        );

    \led7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5839\,
            PADOUT => \N__5838\,
            PADIN => \N__5837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3273\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5830\,
            DIN => \N__5829\,
            DOUT => \N__5828\,
            PACKAGEPIN => lcol1_wire
        );

    \lcol1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5830\,
            PADOUT => \N__5829\,
            PADIN => \N__5828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3768\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1401\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5807\
        );

    \I__1400\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5804\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__5807\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__5804\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1397\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5790\
        );

    \I__1396\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5790\
        );

    \I__1395\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5790\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__5790\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__5787\,
            I => \N__5784\
        );

    \I__1392\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__5781\,
            I => \arse.divseven.doutZ0Z_0\
        );

    \I__1390\ : IoInMux
    port map (
            O => \N__5778\,
            I => \N__5775\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__5775\,
            I => \arse.divseven.dout_i_0\
        );

    \I__1388\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5769\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5764\
        );

    \I__1386\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5761\
        );

    \I__1385\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5758\
        );

    \I__1384\ : Odrv12
    port map (
            O => \N__5764\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__5761\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__5758\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1381\ : ClkMux
    port map (
            O => \N__5751\,
            I => \N__5709\
        );

    \I__1380\ : ClkMux
    port map (
            O => \N__5750\,
            I => \N__5709\
        );

    \I__1379\ : ClkMux
    port map (
            O => \N__5749\,
            I => \N__5709\
        );

    \I__1378\ : ClkMux
    port map (
            O => \N__5748\,
            I => \N__5709\
        );

    \I__1377\ : ClkMux
    port map (
            O => \N__5747\,
            I => \N__5709\
        );

    \I__1376\ : ClkMux
    port map (
            O => \N__5746\,
            I => \N__5709\
        );

    \I__1375\ : ClkMux
    port map (
            O => \N__5745\,
            I => \N__5709\
        );

    \I__1374\ : ClkMux
    port map (
            O => \N__5744\,
            I => \N__5709\
        );

    \I__1373\ : ClkMux
    port map (
            O => \N__5743\,
            I => \N__5709\
        );

    \I__1372\ : ClkMux
    port map (
            O => \N__5742\,
            I => \N__5709\
        );

    \I__1371\ : ClkMux
    port map (
            O => \N__5741\,
            I => \N__5709\
        );

    \I__1370\ : ClkMux
    port map (
            O => \N__5740\,
            I => \N__5709\
        );

    \I__1369\ : ClkMux
    port map (
            O => \N__5739\,
            I => \N__5709\
        );

    \I__1368\ : ClkMux
    port map (
            O => \N__5738\,
            I => \N__5709\
        );

    \I__1367\ : GlobalMux
    port map (
            O => \N__5709\,
            I => \N__5706\
        );

    \I__1366\ : gio2CtrlBuf
    port map (
            O => \N__5706\,
            I => \PLLOUTCORE_g\
        );

    \I__1365\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__5700\,
            I => \arse.divseven.doutZ0Z_1\
        );

    \I__1363\ : IoInMux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__5694\,
            I => \arse.divseven.dout_i_1\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__5691\,
            I => \N__5685\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5678\
        );

    \I__1359\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5678\
        );

    \I__1358\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5675\
        );

    \I__1357\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5672\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \N__5669\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__5683\,
            I => \N__5666\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__5678\,
            I => \N__5659\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5659\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5659\
        );

    \I__1351\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5656\
        );

    \I__1350\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5653\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__5659\,
            I => \N__5650\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__5656\,
            I => \N__5646\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5643\
        );

    \I__1346\ : Span4Mux_h
    port map (
            O => \N__5650\,
            I => \N__5640\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__5649\,
            I => \N__5637\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__5646\,
            I => \N__5634\
        );

    \I__1343\ : Span12Mux_v
    port map (
            O => \N__5643\,
            I => \N__5631\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__5640\,
            I => \N__5628\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5625\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__5634\,
            I => \delayConstantZ0Z_2\
        );

    \I__1339\ : Odrv12
    port map (
            O => \N__5631\,
            I => \delayConstantZ0Z_2\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__5628\,
            I => \delayConstantZ0Z_2\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5625\,
            I => \delayConstantZ0Z_2\
        );

    \I__1336\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5606\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5603\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5594\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5594\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5594\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5594\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5589\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5589\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__5606\,
            I => \N__5583\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5603\,
            I => \N__5580\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5575\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__5589\,
            I => \N__5575\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5572\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5566\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5566\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__5583\,
            I => \N__5563\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__5580\,
            I => \N__5558\
        );

    \I__1319\ : Span4Mux_v
    port map (
            O => \N__5575\,
            I => \N__5558\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5572\,
            I => \N__5555\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__5571\,
            I => \N__5552\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5549\
        );

    \I__1315\ : Span4Mux_h
    port map (
            O => \N__5563\,
            I => \N__5546\
        );

    \I__1314\ : Sp12to4
    port map (
            O => \N__5558\,
            I => \N__5543\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__5555\,
            I => \N__5540\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5537\
        );

    \I__1311\ : Span12Mux_v
    port map (
            O => \N__5549\,
            I => \N__5534\
        );

    \I__1310\ : Sp12to4
    port map (
            O => \N__5546\,
            I => \N__5529\
        );

    \I__1309\ : Span12Mux_h
    port map (
            O => \N__5543\,
            I => \N__5529\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__5540\,
            I => \delayConstantZ0Z_1\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5537\,
            I => \delayConstantZ0Z_1\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__5534\,
            I => \delayConstantZ0Z_1\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__5529\,
            I => \delayConstantZ0Z_1\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5517\,
            I => \N__5509\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5506\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5503\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5496\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5496\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5496\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__5509\,
            I => arse_cpuclkreset
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5506\,
            I => arse_cpuclkreset
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5503\,
            I => arse_cpuclkreset
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5496\,
            I => arse_cpuclkreset
        );

    \I__1293\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5484\,
            I => apusync_c
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__5481\,
            I => \N__5477\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5474\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5471\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5474\,
            I => \N__5464\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5471\,
            I => \N__5464\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5459\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5459\
        );

    \I__1284\ : Span4Mux_h
    port map (
            O => \N__5464\,
            I => \N__5454\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5454\
        );

    \I__1282\ : Span4Mux_v
    port map (
            O => \N__5454\,
            I => \N__5450\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5447\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__5450\,
            I => \arse.apusynclatchedZ0\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5447\,
            I => \arse.apusynclatchedZ0\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5439\,
            I => \arse.diveight.doutZ0Z_0\
        );

    \I__1276\ : IoInMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5433\,
            I => \arse.diveight.dout_i_0\
        );

    \I__1274\ : IoInMux
    port map (
            O => \N__5430\,
            I => \N__5427\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5427\,
            I => \arse.diveight.dout_i_1\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5421\,
            I => \N__5417\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5414\
        );

    \I__1269\ : Span4Mux_s0_h
    port map (
            O => \N__5417\,
            I => \N__5408\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5408\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5405\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__5408\,
            I => \N__5402\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5399\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__5402\,
            I => \N__5396\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__5399\,
            I => \N__5393\
        );

    \I__1262\ : Sp12to4
    port map (
            O => \N__5396\,
            I => \N__5388\
        );

    \I__1261\ : Sp12to4
    port map (
            O => \N__5393\,
            I => \N__5388\
        );

    \I__1260\ : Span12Mux_h
    port map (
            O => \N__5388\,
            I => \N__5384\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5381\
        );

    \I__1258\ : Odrv12
    port map (
            O => \N__5384\,
            I => debouncedconsolereset
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5381\,
            I => debouncedconsolereset
        );

    \I__1256\ : IoInMux
    port map (
            O => \N__5376\,
            I => \N__5373\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5373\,
            I => \arse.apuresetoutregZ0\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5365\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5360\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5360\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5365\,
            I => arse_diveight_counter_1
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5360\,
            I => arse_diveight_counter_1
        );

    \I__1249\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5349\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5346\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5341\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5341\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5349\,
            I => arse_diveight_counter_0
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5346\,
            I => arse_diveight_counter_0
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5341\,
            I => arse_diveight_counter_0
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5328\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5328\,
            I => \N__5322\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5319\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__5326\,
            I => \N__5316\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__5325\,
            I => \N__5308\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__5322\,
            I => \N__5303\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5319\,
            I => \N__5303\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5300\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__5315\,
            I => \N__5297\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__5314\,
            I => \N__5294\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__5313\,
            I => \N__5290\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__5312\,
            I => \N__5287\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__5311\,
            I => \N__5284\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5279\
        );

    \I__1227\ : Span4Mux_h
    port map (
            O => \N__5303\,
            I => \N__5274\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5274\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5271\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5264\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5264\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5264\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5259\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5284\,
            I => \N__5259\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5256\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5253\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5279\,
            I => \N__5250\
        );

    \I__1216\ : Span4Mux_h
    port map (
            O => \N__5274\,
            I => \N__5247\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5271\,
            I => \N__5240\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5264\,
            I => \N__5240\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5259\,
            I => \N__5240\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5256\,
            I => \N__5235\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5253\,
            I => \N__5228\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__5250\,
            I => \N__5228\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__5247\,
            I => \N__5228\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__5240\,
            I => \N__5225\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5220\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5220\
        );

    \I__1205\ : Span4Mux_h
    port map (
            O => \N__5235\,
            I => \N__5217\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__5228\,
            I => \delayConstantZ0Z_0\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__5225\,
            I => \delayConstantZ0Z_0\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5220\,
            I => \delayConstantZ0Z_0\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__5217\,
            I => \delayConstantZ0Z_0\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5203\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5200\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5197\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5203\,
            I => arse_diveight_counter_2
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5200\,
            I => arse_diveight_counter_2
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5197\,
            I => arse_diveight_counter_2
        );

    \I__1194\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5187\,
            I => \arse.diveight.doutZ0Z_1\
        );

    \I__1192\ : SRMux
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5181\,
            I => \N__5178\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__5178\,
            I => \arse.diveight.cpuclkreset_i\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__5175\,
            I => \arse.m8_2_cascade_\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5167\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5162\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5162\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5167\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5162\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__5157\,
            I => \N__5152\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5149\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5144\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5144\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5149\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5144\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__5139\,
            I => \N__5135\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5131\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5126\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5126\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5131\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5126\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5116\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5111\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5111\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5116\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5111\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__5106\,
            I => \arse.m12_2_cascade_\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5098\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5095\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5092\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5098\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5095\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5092\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5082\,
            I => \arse.cpuresetoutreg_1_sqmuxa\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5075\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5072\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5075\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5072\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5063\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5060\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5063\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5060\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5051\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5048\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5051\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5048\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5037\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5037\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5037\,
            I => \arse.m4_e_2\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5031\,
            I => \arse.cpuclkreset_1_sqmuxa\
        );

    \I__1140\ : SRMux
    port map (
            O => \N__5028\,
            I => \N__5023\
        );

    \I__1139\ : SRMux
    port map (
            O => \N__5027\,
            I => \N__5020\
        );

    \I__1138\ : SRMux
    port map (
            O => \N__5026\,
            I => \N__5017\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5023\,
            I => \N__5014\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5020\,
            I => \N__5011\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__5008\
        );

    \I__1134\ : Span4Mux_v
    port map (
            O => \N__5014\,
            I => \N__5005\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__5011\,
            I => debouncedconsolereset_i
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__5008\,
            I => debouncedconsolereset_i
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__5005\,
            I => debouncedconsolereset_i
        );

    \I__1130\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4991\
        );

    \I__1129\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4987\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4984\
        );

    \I__1127\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4981\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__4994\,
            I => \N__4978\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4975\
        );

    \I__1124\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4972\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__4987\,
            I => \N__4968\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__4984\,
            I => \N__4965\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__4981\,
            I => \N__4962\
        );

    \I__1120\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4959\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__4975\,
            I => \N__4956\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4953\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__4971\,
            I => \N__4950\
        );

    \I__1116\ : Sp12to4
    port map (
            O => \N__4968\,
            I => \N__4941\
        );

    \I__1115\ : Sp12to4
    port map (
            O => \N__4965\,
            I => \N__4941\
        );

    \I__1114\ : Sp12to4
    port map (
            O => \N__4962\,
            I => \N__4941\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__4959\,
            I => \N__4941\
        );

    \I__1112\ : Span4Mux_h
    port map (
            O => \N__4956\,
            I => \N__4938\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__4953\,
            I => \N__4935\
        );

    \I__1110\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4932\
        );

    \I__1109\ : Span12Mux_v
    port map (
            O => \N__4941\,
            I => \N__4929\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__4938\,
            I => \N__4926\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__4935\,
            I => \delayConstantZ0Z_3\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__4932\,
            I => \delayConstantZ0Z_3\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__4929\,
            I => \delayConstantZ0Z_3\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__4926\,
            I => \delayConstantZ0Z_3\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__4917\,
            I => \arse_diveight_N_123_0_cascade_\
        );

    \I__1102\ : InMux
    port map (
            O => \N__4914\,
            I => \arse.un1_cpuresetcount_1_cry_1\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4911\,
            I => \arse.un1_cpuresetcount_1_cry_2\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4908\,
            I => \arse.un1_cpuresetcount_1_cry_3\
        );

    \I__1099\ : InMux
    port map (
            O => \N__4905\,
            I => \arse.un1_cpuresetcount_1_cry_4\
        );

    \I__1098\ : InMux
    port map (
            O => \N__4902\,
            I => \arse.un1_cpuresetcount_1_cry_5\
        );

    \I__1097\ : InMux
    port map (
            O => \N__4899\,
            I => \arse.un1_cpuresetcount_1_cry_6\
        );

    \I__1096\ : IoInMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__4893\,
            I => \N__4889\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4886\
        );

    \I__1093\ : Span12Mux_s2_h
    port map (
            O => \N__4889\,
            I => \N__4883\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__4886\,
            I => \arse.cpuresetoutregZ0\
        );

    \I__1091\ : Odrv12
    port map (
            O => \N__4883\,
            I => \arse.cpuresetoutregZ0\
        );

    \I__1090\ : IoInMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__1088\ : Span4Mux_s2_v
    port map (
            O => \N__4872\,
            I => \N__4868\
        );

    \I__1087\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4865\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__4868\,
            I => \N__4860\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__4865\,
            I => \N__4857\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__4864\,
            I => \N__4854\
        );

    \I__1083\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4849\
        );

    \I__1082\ : Span4Mux_h
    port map (
            O => \N__4860\,
            I => \N__4846\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__4857\,
            I => \N__4843\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4838\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4838\
        );

    \I__1078\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4835\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4849\,
            I => \N__4831\
        );

    \I__1076\ : Sp12to4
    port map (
            O => \N__4846\,
            I => \N__4828\
        );

    \I__1075\ : Span12Mux_v
    port map (
            O => \N__4843\,
            I => \N__4825\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__4838\,
            I => \N__4822\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4819\
        );

    \I__1072\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4816\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__4831\,
            I => \N__4813\
        );

    \I__1070\ : Span12Mux_v
    port map (
            O => \N__4828\,
            I => \N__4810\
        );

    \I__1069\ : Span12Mux_h
    port map (
            O => \N__4825\,
            I => \N__4807\
        );

    \I__1068\ : Span12Mux_h
    port map (
            O => \N__4822\,
            I => \N__4802\
        );

    \I__1067\ : Span12Mux_v
    port map (
            O => \N__4819\,
            I => \N__4802\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__4816\,
            I => \N__4797\
        );

    \I__1065\ : Sp12to4
    port map (
            O => \N__4813\,
            I => \N__4797\
        );

    \I__1064\ : Span12Mux_v
    port map (
            O => \N__4810\,
            I => \N__4792\
        );

    \I__1063\ : Span12Mux_h
    port map (
            O => \N__4807\,
            I => \N__4792\
        );

    \I__1062\ : Span12Mux_v
    port map (
            O => \N__4802\,
            I => \N__4789\
        );

    \I__1061\ : Span12Mux_h
    port map (
            O => \N__4797\,
            I => \N__4786\
        );

    \I__1060\ : Odrv12
    port map (
            O => \N__4792\,
            I => masterreset_c
        );

    \I__1059\ : Odrv12
    port map (
            O => \N__4789\,
            I => masterreset_c
        );

    \I__1058\ : Odrv12
    port map (
            O => \N__4786\,
            I => masterreset_c
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__4779\,
            I => \delayConstant17_i_cascade_\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4773\,
            I => \un1_delayConstant_cry_0_c_RNOZ0\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__4767\,
            I => \olddn_RNIM5BH1Z0Z_4\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4761\,
            I => \olddn_RNIM5BHZ0Z1\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4755\,
            I => \N__4752\
        );

    \I__1048\ : Span12Mux_v
    port map (
            O => \N__4752\,
            I => \N__4742\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4739\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4726\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4726\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4726\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4726\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4726\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4726\
        );

    \I__1040\ : Odrv12
    port map (
            O => \N__4742\,
            I => \olddn_RNIEENHZ0\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4739\,
            I => \olddn_RNIEENHZ0\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4726\,
            I => \olddn_RNIEENHZ0\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4716\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__1035\ : Span4Mux_h
    port map (
            O => \N__4713\,
            I => \N__4707\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__4712\,
            I => \N__4703\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__4711\,
            I => \N__4699\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__4710\,
            I => \N__4696\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__4707\,
            I => \N__4691\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4688\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4677\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4677\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4677\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4677\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4677\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4674\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__4691\,
            I => \delayConstant17_i\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4688\,
            I => \delayConstant17_i\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4677\,
            I => \delayConstant17_i\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4674\,
            I => \delayConstant17_i\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4662\,
            I => \olddn_RNIM5BH1Z0Z_2\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4656\,
            I => \oldupZ0\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4649\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__4652\,
            I => \N__4646\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__1011\ : Span12Mux_s9_h
    port map (
            O => \N__4643\,
            I => \N__4637\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4640\,
            I => \debounceup.counter19\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__4637\,
            I => \debounceup.counter19\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__1006\ : Span4Mux_v
    port map (
            O => \N__4626\,
            I => \N__4623\
        );

    \I__1005\ : Sp12to4
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__1004\ : Span12Mux_s6_h
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__1003\ : Odrv12
    port map (
            O => \N__4617\,
            I => delup_c
        );

    \I__1002\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4610\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4607\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4588\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4585\
        );

    \I__998\ : CEMux
    port map (
            O => \N__4606\,
            I => \N__4548\
        );

    \I__997\ : CEMux
    port map (
            O => \N__4605\,
            I => \N__4548\
        );

    \I__996\ : CEMux
    port map (
            O => \N__4604\,
            I => \N__4548\
        );

    \I__995\ : CEMux
    port map (
            O => \N__4603\,
            I => \N__4548\
        );

    \I__994\ : CEMux
    port map (
            O => \N__4602\,
            I => \N__4548\
        );

    \I__993\ : CEMux
    port map (
            O => \N__4601\,
            I => \N__4548\
        );

    \I__992\ : CEMux
    port map (
            O => \N__4600\,
            I => \N__4548\
        );

    \I__991\ : CEMux
    port map (
            O => \N__4599\,
            I => \N__4548\
        );

    \I__990\ : CEMux
    port map (
            O => \N__4598\,
            I => \N__4548\
        );

    \I__989\ : CEMux
    port map (
            O => \N__4597\,
            I => \N__4548\
        );

    \I__988\ : CEMux
    port map (
            O => \N__4596\,
            I => \N__4548\
        );

    \I__987\ : CEMux
    port map (
            O => \N__4595\,
            I => \N__4548\
        );

    \I__986\ : CEMux
    port map (
            O => \N__4594\,
            I => \N__4548\
        );

    \I__985\ : CEMux
    port map (
            O => \N__4593\,
            I => \N__4548\
        );

    \I__984\ : CEMux
    port map (
            O => \N__4592\,
            I => \N__4548\
        );

    \I__983\ : CEMux
    port map (
            O => \N__4591\,
            I => \N__4548\
        );

    \I__982\ : Glb2LocalMux
    port map (
            O => \N__4588\,
            I => \N__4548\
        );

    \I__981\ : Glb2LocalMux
    port map (
            O => \N__4585\,
            I => \N__4548\
        );

    \I__980\ : GlobalMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__979\ : gio2CtrlBuf
    port map (
            O => \N__4545\,
            I => \N_111_g\
        );

    \I__978\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4535\
        );

    \I__977\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4535\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__4540\,
            I => \N__4532\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4529\
        );

    \I__974\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4526\
        );

    \I__973\ : Span12Mux_s10_v
    port map (
            O => \N__4529\,
            I => \N__4523\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4526\,
            I => debouncedup
        );

    \I__971\ : Odrv12
    port map (
            O => \N__4523\,
            I => debouncedup
        );

    \I__970\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4515\,
            I => \N__4484\
        );

    \I__968\ : ClkMux
    port map (
            O => \N__4514\,
            I => \N__4425\
        );

    \I__967\ : ClkMux
    port map (
            O => \N__4513\,
            I => \N__4425\
        );

    \I__966\ : ClkMux
    port map (
            O => \N__4512\,
            I => \N__4425\
        );

    \I__965\ : ClkMux
    port map (
            O => \N__4511\,
            I => \N__4425\
        );

    \I__964\ : ClkMux
    port map (
            O => \N__4510\,
            I => \N__4425\
        );

    \I__963\ : ClkMux
    port map (
            O => \N__4509\,
            I => \N__4425\
        );

    \I__962\ : ClkMux
    port map (
            O => \N__4508\,
            I => \N__4425\
        );

    \I__961\ : ClkMux
    port map (
            O => \N__4507\,
            I => \N__4425\
        );

    \I__960\ : ClkMux
    port map (
            O => \N__4506\,
            I => \N__4425\
        );

    \I__959\ : ClkMux
    port map (
            O => \N__4505\,
            I => \N__4425\
        );

    \I__958\ : ClkMux
    port map (
            O => \N__4504\,
            I => \N__4425\
        );

    \I__957\ : ClkMux
    port map (
            O => \N__4503\,
            I => \N__4425\
        );

    \I__956\ : ClkMux
    port map (
            O => \N__4502\,
            I => \N__4425\
        );

    \I__955\ : ClkMux
    port map (
            O => \N__4501\,
            I => \N__4425\
        );

    \I__954\ : ClkMux
    port map (
            O => \N__4500\,
            I => \N__4425\
        );

    \I__953\ : ClkMux
    port map (
            O => \N__4499\,
            I => \N__4425\
        );

    \I__952\ : ClkMux
    port map (
            O => \N__4498\,
            I => \N__4425\
        );

    \I__951\ : ClkMux
    port map (
            O => \N__4497\,
            I => \N__4425\
        );

    \I__950\ : ClkMux
    port map (
            O => \N__4496\,
            I => \N__4425\
        );

    \I__949\ : ClkMux
    port map (
            O => \N__4495\,
            I => \N__4425\
        );

    \I__948\ : ClkMux
    port map (
            O => \N__4494\,
            I => \N__4425\
        );

    \I__947\ : ClkMux
    port map (
            O => \N__4493\,
            I => \N__4425\
        );

    \I__946\ : ClkMux
    port map (
            O => \N__4492\,
            I => \N__4425\
        );

    \I__945\ : ClkMux
    port map (
            O => \N__4491\,
            I => \N__4425\
        );

    \I__944\ : ClkMux
    port map (
            O => \N__4490\,
            I => \N__4425\
        );

    \I__943\ : ClkMux
    port map (
            O => \N__4489\,
            I => \N__4425\
        );

    \I__942\ : ClkMux
    port map (
            O => \N__4488\,
            I => \N__4425\
        );

    \I__941\ : ClkMux
    port map (
            O => \N__4487\,
            I => \N__4425\
        );

    \I__940\ : Glb2LocalMux
    port map (
            O => \N__4484\,
            I => \N__4425\
        );

    \I__939\ : GlobalMux
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__938\ : gio2CtrlBuf
    port map (
            O => \N__4422\,
            I => \PACKAGEPIN_0_c_g\
        );

    \I__937\ : InMux
    port map (
            O => \N__4419\,
            I => \arse.un1_cpuresetcount_1_cry_0\
        );

    \I__936\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4409\
        );

    \I__935\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4406\
        );

    \I__934\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4400\
        );

    \I__933\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4395\
        );

    \I__932\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4395\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4390\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4390\
        );

    \I__929\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4385\
        );

    \I__928\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4385\
        );

    \I__927\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4381\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4376\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4395\,
            I => \N__4376\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__4390\,
            I => \N__4369\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4385\,
            I => \N__4369\
        );

    \I__922\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4366\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4381\,
            I => \N__4363\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__4376\,
            I => \N__4360\
        );

    \I__919\ : InMux
    port map (
            O => \N__4375\,
            I => \N__4357\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__4374\,
            I => \N__4354\
        );

    \I__917\ : Span4Mux_h
    port map (
            O => \N__4369\,
            I => \N__4351\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4366\,
            I => \N__4342\
        );

    \I__915\ : Sp12to4
    port map (
            O => \N__4363\,
            I => \N__4342\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__4360\,
            I => \N__4342\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4357\,
            I => \N__4342\
        );

    \I__912\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4339\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__4351\,
            I => \N__4336\
        );

    \I__910\ : Span12Mux_v
    port map (
            O => \N__4342\,
            I => \N__4333\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4339\,
            I => \delayConstantZ0Z_4\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__4336\,
            I => \delayConstantZ0Z_4\
        );

    \I__907\ : Odrv12
    port map (
            O => \N__4333\,
            I => \delayConstantZ0Z_4\
        );

    \I__906\ : InMux
    port map (
            O => \N__4326\,
            I => \un1_delayConstant_cry_3\
        );

    \I__905\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4318\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4322\,
            I => \N__4315\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__4321\,
            I => \N__4312\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4318\,
            I => \N__4308\
        );

    \I__901\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4305\
        );

    \I__900\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4300\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__4311\,
            I => \N__4296\
        );

    \I__898\ : Span4Mux_v
    port map (
            O => \N__4308\,
            I => \N__4289\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4289\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__4304\,
            I => \N__4286\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__4303\,
            I => \N__4282\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4300\,
            I => \N__4279\
        );

    \I__893\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4274\
        );

    \I__892\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4274\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__4295\,
            I => \N__4271\
        );

    \I__890\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4268\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__4289\,
            I => \N__4265\
        );

    \I__888\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4260\
        );

    \I__887\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4260\
        );

    \I__886\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4256\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__4279\,
            I => \N__4253\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4274\,
            I => \N__4250\
        );

    \I__883\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4247\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4244\
        );

    \I__881\ : Span4Mux_h
    port map (
            O => \N__4265\,
            I => \N__4239\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4260\,
            I => \N__4239\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4259\,
            I => \N__4236\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4256\,
            I => \N__4231\
        );

    \I__877\ : Sp12to4
    port map (
            O => \N__4253\,
            I => \N__4231\
        );

    \I__876\ : Sp12to4
    port map (
            O => \N__4250\,
            I => \N__4226\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4247\,
            I => \N__4226\
        );

    \I__874\ : Span4Mux_v
    port map (
            O => \N__4244\,
            I => \N__4223\
        );

    \I__873\ : Span4Mux_h
    port map (
            O => \N__4239\,
            I => \N__4220\
        );

    \I__872\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4217\
        );

    \I__871\ : Span12Mux_h
    port map (
            O => \N__4231\,
            I => \N__4214\
        );

    \I__870\ : Span12Mux_v
    port map (
            O => \N__4226\,
            I => \N__4211\
        );

    \I__869\ : Span4Mux_h
    port map (
            O => \N__4223\,
            I => \N__4206\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__4220\,
            I => \N__4206\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4217\,
            I => \delayConstantZ0Z_5\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__4214\,
            I => \delayConstantZ0Z_5\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__4211\,
            I => \delayConstantZ0Z_5\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__4206\,
            I => \delayConstantZ0Z_5\
        );

    \I__863\ : InMux
    port map (
            O => \N__4197\,
            I => \un1_delayConstant_cry_4\
        );

    \I__862\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4191\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4191\,
            I => \N__4187\
        );

    \I__860\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4182\
        );

    \I__859\ : Span4Mux_h
    port map (
            O => \N__4187\,
            I => \N__4178\
        );

    \I__858\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4175\
        );

    \I__857\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4172\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4182\,
            I => \N__4168\
        );

    \I__855\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4165\
        );

    \I__854\ : Span4Mux_h
    port map (
            O => \N__4178\,
            I => \N__4160\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4175\,
            I => \N__4160\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4172\,
            I => \N__4157\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \N__4154\
        );

    \I__850\ : Sp12to4
    port map (
            O => \N__4168\,
            I => \N__4149\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4149\
        );

    \I__848\ : Span4Mux_h
    port map (
            O => \N__4160\,
            I => \N__4146\
        );

    \I__847\ : Span12Mux_h
    port map (
            O => \N__4157\,
            I => \N__4143\
        );

    \I__846\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4140\
        );

    \I__845\ : Span12Mux_v
    port map (
            O => \N__4149\,
            I => \N__4137\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__4146\,
            I => \N__4134\
        );

    \I__843\ : Odrv12
    port map (
            O => \N__4143\,
            I => \delayConstantZ0Z_6\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4140\,
            I => \delayConstantZ0Z_6\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__4137\,
            I => \delayConstantZ0Z_6\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4134\,
            I => \delayConstantZ0Z_6\
        );

    \I__839\ : InMux
    port map (
            O => \N__4125\,
            I => \un1_delayConstant_cry_5\
        );

    \I__838\ : InMux
    port map (
            O => \N__4122\,
            I => \un1_delayConstant_cry_6\
        );

    \I__837\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4115\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__4118\,
            I => \N__4111\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4115\,
            I => \N__4106\
        );

    \I__834\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4101\
        );

    \I__833\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4101\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__4110\,
            I => \N__4098\
        );

    \I__831\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4095\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__4106\,
            I => \N__4090\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4101\,
            I => \N__4090\
        );

    \I__828\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4086\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4083\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__4090\,
            I => \N__4080\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4089\,
            I => \N__4077\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4086\,
            I => \N__4074\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__4083\,
            I => \N__4069\
        );

    \I__822\ : Span4Mux_h
    port map (
            O => \N__4080\,
            I => \N__4069\
        );

    \I__821\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4066\
        );

    \I__820\ : Span12Mux_h
    port map (
            O => \N__4074\,
            I => \N__4063\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__4069\,
            I => \N__4060\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4066\,
            I => \delayConstantZ0Z_7\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__4063\,
            I => \delayConstantZ0Z_7\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__4060\,
            I => \delayConstantZ0Z_7\
        );

    \I__815\ : SRMux
    port map (
            O => \N__4053\,
            I => \N__4035\
        );

    \I__814\ : SRMux
    port map (
            O => \N__4052\,
            I => \N__4035\
        );

    \I__813\ : SRMux
    port map (
            O => \N__4051\,
            I => \N__4035\
        );

    \I__812\ : SRMux
    port map (
            O => \N__4050\,
            I => \N__4035\
        );

    \I__811\ : SRMux
    port map (
            O => \N__4049\,
            I => \N__4035\
        );

    \I__810\ : SRMux
    port map (
            O => \N__4048\,
            I => \N__4035\
        );

    \I__809\ : GlobalMux
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__808\ : gio2CtrlBuf
    port map (
            O => \N__4032\,
            I => masterreset_c_i_g
        );

    \I__807\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4026\,
            I => \olddnZ0\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__804\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4015\
        );

    \I__803\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4010\
        );

    \I__802\ : InMux
    port map (
            O => \N__4018\,
            I => \N__4010\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4015\,
            I => debounceddn
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4010\,
            I => debounceddn
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__4005\,
            I => \olddn_RNIEENHZ0_cascade_\
        );

    \I__798\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3999\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__3999\,
            I => \olddn_RNIM5BH1Z0Z_0\
        );

    \I__796\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3993\,
            I => \olddn_RNIM5BH1Z0Z_3\
        );

    \I__794\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3987\,
            I => \olddn_RNIM5BH1Z0Z_1\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__3984\,
            I => \N__3981\
        );

    \I__791\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3976\
        );

    \I__790\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3973\
        );

    \I__789\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3970\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__3976\,
            I => \N__3965\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__3973\,
            I => \N__3965\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3970\,
            I => \debouncedn.counter19_2\
        );

    \I__785\ : Odrv4
    port map (
            O => \N__3965\,
            I => \debouncedn.counter19_2\
        );

    \I__784\ : InMux
    port map (
            O => \N__3960\,
            I => \debouncedn.un3_counter_1_cry_3\
        );

    \I__783\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3951\
        );

    \I__782\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3948\
        );

    \I__781\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3945\
        );

    \I__780\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3942\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3951\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3948\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__3945\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3942\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__775\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3927\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__3932\,
            I => \N__3924\
        );

    \I__773\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3921\
        );

    \I__772\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3918\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3927\,
            I => \N__3915\
        );

    \I__770\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3912\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__3921\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3918\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__3915\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3912\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__765\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3899\
        );

    \I__764\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3895\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3899\,
            I => \N__3892\
        );

    \I__762\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3889\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3895\,
            I => \debouncedn.counterZ0Z_1\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3892\,
            I => \debouncedn.counterZ0Z_1\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3889\,
            I => \debouncedn.counterZ0Z_1\
        );

    \I__758\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3879\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3879\,
            I => \N__3875\
        );

    \I__756\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3872\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__3875\,
            I => \N__3869\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3872\,
            I => \debouncedn.counter19\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__3869\,
            I => \debouncedn.counter19\
        );

    \I__752\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__749\ : Span4Mux_h
    port map (
            O => \N__3855\,
            I => \N__3852\
        );

    \I__748\ : Sp12to4
    port map (
            O => \N__3852\,
            I => \N__3849\
        );

    \I__747\ : Span12Mux_h
    port map (
            O => \N__3849\,
            I => \N__3846\
        );

    \I__746\ : Span12Mux_v
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__745\ : Odrv12
    port map (
            O => \N__3843\,
            I => deldn_c
        );

    \I__744\ : IoInMux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3837\,
            I => \N__3833\
        );

    \I__742\ : IoInMux
    port map (
            O => \N__3836\,
            I => \N__3829\
        );

    \I__741\ : IoSpan4Mux
    port map (
            O => \N__3833\,
            I => \N__3826\
        );

    \I__740\ : IoInMux
    port map (
            O => \N__3832\,
            I => \N__3823\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3829\,
            I => \N__3820\
        );

    \I__738\ : IoSpan4Mux
    port map (
            O => \N__3826\,
            I => \N__3814\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3823\,
            I => \N__3814\
        );

    \I__736\ : IoSpan4Mux
    port map (
            O => \N__3820\,
            I => \N__3811\
        );

    \I__735\ : IoInMux
    port map (
            O => \N__3819\,
            I => \N__3808\
        );

    \I__734\ : IoSpan4Mux
    port map (
            O => \N__3814\,
            I => \N__3805\
        );

    \I__733\ : IoSpan4Mux
    port map (
            O => \N__3811\,
            I => \N__3800\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3808\,
            I => \N__3800\
        );

    \I__731\ : Span4Mux_s0_h
    port map (
            O => \N__3805\,
            I => \N__3797\
        );

    \I__730\ : IoSpan4Mux
    port map (
            O => \N__3800\,
            I => \N__3794\
        );

    \I__729\ : Sp12to4
    port map (
            O => \N__3797\,
            I => \N__3791\
        );

    \I__728\ : Span4Mux_s3_v
    port map (
            O => \N__3794\,
            I => \N__3788\
        );

    \I__727\ : Span12Mux_v
    port map (
            O => \N__3791\,
            I => \N__3785\
        );

    \I__726\ : Span4Mux_v
    port map (
            O => \N__3788\,
            I => \N__3782\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__3785\,
            I => \CONSTANT_ONE_NET\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__3782\,
            I => \CONSTANT_ONE_NET\
        );

    \I__723\ : InMux
    port map (
            O => \N__3777\,
            I => \un1_delayConstant_cry_0\
        );

    \I__722\ : InMux
    port map (
            O => \N__3774\,
            I => \un1_delayConstant_cry_1\
        );

    \I__721\ : InMux
    port map (
            O => \N__3771\,
            I => \un1_delayConstant_cry_2\
        );

    \I__720\ : IoInMux
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__718\ : Span4Mux_s2_v
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__717\ : Span4Mux_h
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__3756\,
            I => lcol1_c
        );

    \I__715\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3749\
        );

    \I__714\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3746\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3749\,
            I => \N__3740\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3746\,
            I => \N__3740\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__3745\,
            I => \N__3733\
        );

    \I__710\ : Span4Mux_v
    port map (
            O => \N__3740\,
            I => \N__3729\
        );

    \I__709\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3726\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__3738\,
            I => \N__3722\
        );

    \I__707\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3716\
        );

    \I__706\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3711\
        );

    \I__705\ : InMux
    port map (
            O => \N__3733\,
            I => \N__3711\
        );

    \I__704\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3706\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__3729\,
            I => \N__3701\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3726\,
            I => \N__3701\
        );

    \I__701\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3698\
        );

    \I__700\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3693\
        );

    \I__699\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3693\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3720\,
            I => \N__3688\
        );

    \I__697\ : InMux
    port map (
            O => \N__3719\,
            I => \N__3683\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3716\,
            I => \N__3678\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3711\,
            I => \N__3678\
        );

    \I__694\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3673\
        );

    \I__693\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3673\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3706\,
            I => \N__3667\
        );

    \I__691\ : Span12Mux_h
    port map (
            O => \N__3701\,
            I => \N__3667\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3698\,
            I => \N__3661\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3693\,
            I => \N__3661\
        );

    \I__688\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3654\
        );

    \I__687\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3645\
        );

    \I__686\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3645\
        );

    \I__685\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3645\
        );

    \I__684\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3645\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3683\,
            I => \N__3638\
        );

    \I__682\ : Span4Mux_v
    port map (
            O => \N__3678\,
            I => \N__3638\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3673\,
            I => \N__3638\
        );

    \I__680\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3635\
        );

    \I__679\ : Span12Mux_v
    port map (
            O => \N__3667\,
            I => \N__3632\
        );

    \I__678\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3629\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__3661\,
            I => \N__3626\
        );

    \I__676\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3621\
        );

    \I__675\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3621\
        );

    \I__674\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3616\
        );

    \I__673\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3616\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3654\,
            I => \N__3613\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3645\,
            I => \N__3608\
        );

    \I__670\ : Span4Mux_h
    port map (
            O => \N__3638\,
            I => \N__3608\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3635\,
            I => \colZ0Z_1\
        );

    \I__668\ : Odrv12
    port map (
            O => \N__3632\,
            I => \colZ0Z_1\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3629\,
            I => \colZ0Z_1\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__3626\,
            I => \colZ0Z_1\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3621\,
            I => \colZ0Z_1\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3616\,
            I => \colZ0Z_1\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__3613\,
            I => \colZ0Z_1\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__3608\,
            I => \colZ0Z_1\
        );

    \I__661\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3588\,
            I => \N__3583\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__3587\,
            I => \N__3576\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__3586\,
            I => \N__3573\
        );

    \I__657\ : Span4Mux_h
    port map (
            O => \N__3583\,
            I => \N__3568\
        );

    \I__656\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3565\
        );

    \I__655\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3562\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__3580\,
            I => \N__3549\
        );

    \I__653\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3546\
        );

    \I__652\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3541\
        );

    \I__651\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3541\
        );

    \I__650\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3538\
        );

    \I__649\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3535\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__3568\,
            I => \N__3532\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3565\,
            I => \N__3529\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3562\,
            I => \N__3526\
        );

    \I__645\ : InMux
    port map (
            O => \N__3561\,
            I => \N__3517\
        );

    \I__644\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3517\
        );

    \I__643\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3517\
        );

    \I__642\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3517\
        );

    \I__641\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3514\
        );

    \I__640\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3509\
        );

    \I__639\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3509\
        );

    \I__638\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3505\
        );

    \I__637\ : InMux
    port map (
            O => \N__3553\,
            I => \N__3500\
        );

    \I__636\ : InMux
    port map (
            O => \N__3552\,
            I => \N__3500\
        );

    \I__635\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3497\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3492\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3541\,
            I => \N__3492\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3538\,
            I => \N__3489\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3535\,
            I => \N__3479\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__3532\,
            I => \N__3479\
        );

    \I__629\ : Span12Mux_h
    port map (
            O => \N__3529\,
            I => \N__3479\
        );

    \I__628\ : Sp12to4
    port map (
            O => \N__3526\,
            I => \N__3479\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3517\,
            I => \N__3469\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3514\,
            I => \N__3469\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3509\,
            I => \N__3466\
        );

    \I__624\ : InMux
    port map (
            O => \N__3508\,
            I => \N__3463\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3505\,
            I => \N__3458\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3500\,
            I => \N__3458\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3497\,
            I => \N__3453\
        );

    \I__620\ : Span4Mux_h
    port map (
            O => \N__3492\,
            I => \N__3453\
        );

    \I__619\ : Span4Mux_h
    port map (
            O => \N__3489\,
            I => \N__3450\
        );

    \I__618\ : InMux
    port map (
            O => \N__3488\,
            I => \N__3447\
        );

    \I__617\ : Span12Mux_v
    port map (
            O => \N__3479\,
            I => \N__3444\
        );

    \I__616\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3437\
        );

    \I__615\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3437\
        );

    \I__614\ : InMux
    port map (
            O => \N__3476\,
            I => \N__3437\
        );

    \I__613\ : InMux
    port map (
            O => \N__3475\,
            I => \N__3432\
        );

    \I__612\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3432\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__3469\,
            I => \N__3427\
        );

    \I__610\ : Span4Mux_h
    port map (
            O => \N__3466\,
            I => \N__3427\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3463\,
            I => \N__3420\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__3458\,
            I => \N__3420\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__3453\,
            I => \N__3420\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__3450\,
            I => \colZ0Z_0\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3447\,
            I => \colZ0Z_0\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__3444\,
            I => \colZ0Z_0\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3437\,
            I => \colZ0Z_0\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3432\,
            I => \colZ0Z_0\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__3427\,
            I => \colZ0Z_0\
        );

    \I__600\ : Odrv4
    port map (
            O => \N__3420\,
            I => \colZ0Z_0\
        );

    \I__599\ : IoInMux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3402\,
            I => \N__3399\
        );

    \I__597\ : IoSpan4Mux
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__3396\,
            I => lcol2_c
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__3393\,
            I => \debouncedn.counter19_2_cascade_\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__3390\,
            I => \debouncedn.counter19_cascade_\
        );

    \I__593\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3383\
        );

    \I__592\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3380\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3383\,
            I => \debouncedn.counterZ0Z_2\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3380\,
            I => \debouncedn.counterZ0Z_2\
        );

    \I__589\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3372\,
            I => \debouncedn.counter_RNO_0_1_2\
        );

    \I__587\ : InMux
    port map (
            O => \N__3369\,
            I => \debouncedn.un3_counter_1_cry_1\
        );

    \I__586\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3362\
        );

    \I__585\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3359\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3362\,
            I => \debouncedn.counterZ0Z_3\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3359\,
            I => \debouncedn.counterZ0Z_3\
        );

    \I__582\ : InMux
    port map (
            O => \N__3354\,
            I => \debouncedn.un3_counter_1_cry_2\
        );

    \I__581\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3348\,
            I => \N__3344\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3347\,
            I => \N__3339\
        );

    \I__578\ : Span12Mux_v
    port map (
            O => \N__3344\,
            I => \N__3336\
        );

    \I__577\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3331\
        );

    \I__576\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3331\
        );

    \I__575\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3328\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__3336\,
            I => \debounceup.counterZ0Z_0\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3331\,
            I => \debounceup.counterZ0Z_0\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3328\,
            I => \debounceup.counterZ0Z_0\
        );

    \I__571\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3317\
        );

    \I__570\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3314\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3317\,
            I => \N__3308\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3314\,
            I => \N__3308\
        );

    \I__567\ : InMux
    port map (
            O => \N__3313\,
            I => \N__3305\
        );

    \I__566\ : Span4Mux_v
    port map (
            O => \N__3308\,
            I => \N__3302\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3305\,
            I => \N__3297\
        );

    \I__564\ : Span4Mux_h
    port map (
            O => \N__3302\,
            I => \N__3297\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__3297\,
            I => \debounceup.counterZ0Z_1\
        );

    \I__562\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3291\,
            I => \dig2.m49_bm\
        );

    \I__560\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3285\,
            I => \dig2.m49_am\
        );

    \I__558\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3279\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3279\,
            I => \dig2.m33_am\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__3276\,
            I => \dig2.m33_bm_cascade_\
        );

    \I__555\ : IoInMux
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3270\,
            I => \N__3267\
        );

    \I__553\ : Span12Mux_s4_v
    port map (
            O => \N__3267\,
            I => \N__3264\
        );

    \I__552\ : Span12Mux_v
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__551\ : Span12Mux_h
    port map (
            O => \N__3261\,
            I => \N__3258\
        );

    \I__550\ : Odrv12
    port map (
            O => \N__3258\,
            I => leds_1_i_2
        );

    \I__549\ : CascadeMux
    port map (
            O => \N__3255\,
            I => \dig2.N_25_cascade_\
        );

    \I__548\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3249\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3249\,
            I => \dig2.leds_17_i_0_ns_1_2\
        );

    \I__546\ : InMux
    port map (
            O => \N__3246\,
            I => \N__3243\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3243\,
            I => \dig2.i2_mux\
        );

    \I__544\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3237\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3237\,
            I => \debounceconsolereset.counter_RNO_0Z0Z_2\
        );

    \I__542\ : InMux
    port map (
            O => \N__3234\,
            I => \debounceconsolereset.un3_counter_1_cry_1\
        );

    \I__541\ : InMux
    port map (
            O => \N__3231\,
            I => \debounceconsolereset.un3_counter_1_cry_2\
        );

    \I__540\ : InMux
    port map (
            O => \N__3228\,
            I => \debounceconsolereset.un3_counter_1_cry_3\
        );

    \I__539\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3221\
        );

    \I__538\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3218\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3221\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3218\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__535\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3209\
        );

    \I__534\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3206\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3209\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3206\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__3201\,
            I => \N__3197\
        );

    \I__530\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3193\
        );

    \I__529\ : InMux
    port map (
            O => \N__3197\,
            I => \N__3188\
        );

    \I__528\ : InMux
    port map (
            O => \N__3196\,
            I => \N__3188\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3193\,
            I => \debounceconsolereset.counter19_2\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3188\,
            I => \debounceconsolereset.counter19_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3175\
        );

    \I__524\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3175\
        );

    \I__523\ : InMux
    port map (
            O => \N__3181\,
            I => \N__3172\
        );

    \I__522\ : InMux
    port map (
            O => \N__3180\,
            I => \N__3169\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3175\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3172\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3169\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__3162\,
            I => \N__3158\
        );

    \I__517\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3154\
        );

    \I__516\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3151\
        );

    \I__515\ : InMux
    port map (
            O => \N__3157\,
            I => \N__3148\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3154\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3151\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3148\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3141\,
            I => \debounceconsolereset.counter19_2_cascade_\
        );

    \I__510\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3130\
        );

    \I__509\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3130\
        );

    \I__508\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3127\
        );

    \I__507\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3124\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3130\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3127\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3124\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__3117\,
            I => \N__3114\
        );

    \I__502\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3109\
        );

    \I__501\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3106\
        );

    \I__500\ : InMux
    port map (
            O => \N__3112\,
            I => \N__3103\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3109\,
            I => \debounceconsolereset.counter19\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3106\,
            I => \debounceconsolereset.counter19\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3103\,
            I => \debounceconsolereset.counter19\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3096\,
            I => \N__3092\
        );

    \I__495\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3088\
        );

    \I__494\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3083\
        );

    \I__493\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3080\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3088\,
            I => \N__3077\
        );

    \I__491\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3074\
        );

    \I__490\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3071\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3083\,
            I => \N__3068\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3080\,
            I => col_1_1
        );

    \I__487\ : Odrv4
    port map (
            O => \N__3077\,
            I => col_1_1
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3074\,
            I => col_1_1
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3071\,
            I => col_1_1
        );

    \I__484\ : Odrv12
    port map (
            O => \N__3068\,
            I => col_1_1
        );

    \I__483\ : InMux
    port map (
            O => \N__3057\,
            I => \N__3054\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3054\,
            I => \N__3051\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__3051\,
            I => \dig2.m54_bm\
        );

    \I__480\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3045\,
            I => \N__3042\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__3042\,
            I => \dig2.leds_17_i_ns_1_1\
        );

    \I__477\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3036\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__475\ : Span12Mux_h
    port map (
            O => \N__3033\,
            I => \N__3030\
        );

    \I__474\ : Span12Mux_v
    port map (
            O => \N__3030\,
            I => \N__3027\
        );

    \I__473\ : Odrv12
    port map (
            O => \N__3027\,
            I => consolereset_c
        );

    \I__472\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3021\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3021\,
            I => \N__3018\
        );

    \I__470\ : Span4Mux_h
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__3015\,
            I => \N__3012\
        );

    \I__468\ : Span12Mux_v
    port map (
            O => \N__3012\,
            I => \N__3009\
        );

    \I__467\ : Span12Mux_v
    port map (
            O => \N__3009\,
            I => \N__3006\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__3006\,
            I => altreset_c
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3003\,
            I => \debounceconsolereset.out_RNOZ0Z_0_cascade_\
        );

    \I__464\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2997\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2997\,
            I => \clock_out_RNIR6ER\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__2994\,
            I => \clock_out_RNIR6ER_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2988\,
            I => \N__2983\
        );

    \I__459\ : InMux
    port map (
            O => \N__2987\,
            I => \N__2978\
        );

    \I__458\ : InMux
    port map (
            O => \N__2986\,
            I => \N__2978\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__2983\,
            I => \N__2958\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2978\,
            I => \N__2958\
        );

    \I__455\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2951\
        );

    \I__454\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2951\
        );

    \I__453\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2951\
        );

    \I__452\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2942\
        );

    \I__451\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2942\
        );

    \I__450\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2942\
        );

    \I__449\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2942\
        );

    \I__448\ : InMux
    port map (
            O => \N__2970\,
            I => \N__2939\
        );

    \I__447\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2936\
        );

    \I__446\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2929\
        );

    \I__445\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2929\
        );

    \I__444\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2929\
        );

    \I__443\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2922\
        );

    \I__442\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2922\
        );

    \I__441\ : InMux
    port map (
            O => \N__2963\,
            I => \N__2922\
        );

    \I__440\ : Span4Mux_h
    port map (
            O => \N__2958\,
            I => \N__2919\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2951\,
            I => arses_counter8
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2942\,
            I => arses_counter8
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2939\,
            I => arses_counter8
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2936\,
            I => arses_counter8
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2929\,
            I => arses_counter8
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2922\,
            I => arses_counter8
        );

    \I__433\ : Odrv4
    port map (
            O => \N__2919\,
            I => arses_counter8
        );

    \I__432\ : InMux
    port map (
            O => \N__2904\,
            I => \N__2900\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__2903\,
            I => \N__2896\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2900\,
            I => \N__2890\
        );

    \I__429\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2887\
        );

    \I__428\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2884\
        );

    \I__427\ : InMux
    port map (
            O => \N__2895\,
            I => \N__2877\
        );

    \I__426\ : InMux
    port map (
            O => \N__2894\,
            I => \N__2877\
        );

    \I__425\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2877\
        );

    \I__424\ : Span4Mux_h
    port map (
            O => \N__2890\,
            I => \N__2874\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2887\,
            I => slowclk
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2884\,
            I => slowclk
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2877\,
            I => slowclk
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2874\,
            I => slowclk
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__418\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2859\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2859\,
            I => \dig2.m54_am\
        );

    \I__416\ : IoInMux
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2853\,
            I => \N__2850\
        );

    \I__414\ : Span12Mux_s4_v
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__413\ : Span12Mux_v
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__412\ : Odrv12
    port map (
            O => \N__2844\,
            I => leds_1_i_0_1
        );

    \I__411\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2838\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2838\,
            I => \dig2.m75_ns_1\
        );

    \I__409\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2832\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2832\,
            I => \dig2.m69_am\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__406\ : InMux
    port map (
            O => \N__2826\,
            I => \N__2823\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2823\,
            I => \dig2.m69_bm\
        );

    \I__404\ : IoInMux
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__402\ : IoSpan4Mux
    port map (
            O => \N__2814\,
            I => \N__2811\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__2808\,
            I => \N__2805\
        );

    \I__399\ : Span12Mux_s6_v
    port map (
            O => \N__2805\,
            I => \N__2802\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__2802\,
            I => leds_1_i_0_2
        );

    \I__397\ : InMux
    port map (
            O => \N__2799\,
            I => \N__2796\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2796\,
            I => \dig2.N_78\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__394\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2787\,
            I => \dig2.N_76\
        );

    \I__392\ : IoInMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__390\ : IoSpan4Mux
    port map (
            O => \N__2778\,
            I => \N__2775\
        );

    \I__389\ : Span4Mux_s2_v
    port map (
            O => \N__2775\,
            I => \N__2772\
        );

    \I__388\ : Span4Mux_h
    port map (
            O => \N__2772\,
            I => \N__2769\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__386\ : Span12Mux_v
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__2763\,
            I => leds_1_i_0_3
        );

    \I__384\ : CascadeMux
    port map (
            O => \N__2760\,
            I => \dig2.m39_ns_1_cascade_\
        );

    \I__383\ : InMux
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2754\,
            I => \dig2.N_40\
        );

    \I__381\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2748\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2748\,
            I => \dig2.i3_mux\
        );

    \I__379\ : InMux
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2742\,
            I => \dig2.N_59\
        );

    \I__377\ : InMux
    port map (
            O => \N__2739\,
            I => \N__2736\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2736\,
            I => \dig2.leds_17_i_ns_1_2\
        );

    \I__375\ : InMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2730\,
            I => \dig2.m18_am\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2724\,
            I => \N__2721\
        );

    \I__371\ : IoSpan4Mux
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__370\ : Sp12to4
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__369\ : Span12Mux_v
    port map (
            O => \N__2715\,
            I => \N__2712\
        );

    \I__368\ : Span12Mux_h
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__367\ : Odrv12
    port map (
            O => \N__2709\,
            I => leds_1_i_3
        );

    \I__366\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2703\,
            I => \dig2.m13_bm\
        );

    \I__364\ : InMux
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2697\,
            I => \dig2.N_42\
        );

    \I__362\ : InMux
    port map (
            O => \N__2694\,
            I => \N__2690\
        );

    \I__361\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2690\,
            I => \arses.counterZ0Z_11\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2687\,
            I => \arses.counterZ0Z_11\
        );

    \I__358\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2678\
        );

    \I__357\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2675\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2678\,
            I => \arses.counterZ0Z_10\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2675\,
            I => \arses.counterZ0Z_10\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2670\,
            I => \arses.un1_counterlt11_cascade_\
        );

    \I__353\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2663\
        );

    \I__352\ : InMux
    port map (
            O => \N__2666\,
            I => \N__2660\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2663\,
            I => \arses.counterZ0Z_9\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2660\,
            I => \arses.counterZ0Z_9\
        );

    \I__349\ : InMux
    port map (
            O => \N__2655\,
            I => \N__2651\
        );

    \I__348\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2648\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2651\,
            I => \arses.counterZ0Z_14\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2648\,
            I => \arses.counterZ0Z_14\
        );

    \I__345\ : InMux
    port map (
            O => \N__2643\,
            I => \N__2639\
        );

    \I__344\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2636\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2639\,
            I => \arses.counterZ0Z_13\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2636\,
            I => \arses.counterZ0Z_13\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2631\,
            I => \arses.un1_counterlt13_0_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__2628\,
            I => \N__2624\
        );

    \I__339\ : InMux
    port map (
            O => \N__2627\,
            I => \N__2621\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2624\,
            I => \arses.counterZ0Z_12\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2621\,
            I => \arses.counterZ0Z_12\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__2616\,
            I => \arses_counter8_cascade_\
        );

    \I__335\ : IoInMux
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2610\,
            I => \N__2607\
        );

    \I__333\ : Span4Mux_s2_v
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__2604\,
            I => \N__2601\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__2601\,
            I => \arses.clock_out_RNIR6ERZ0Z_0\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__329\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2592\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2592\,
            I => \N__2587\
        );

    \I__327\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2582\
        );

    \I__326\ : InMux
    port map (
            O => \N__2590\,
            I => \N__2582\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__2587\,
            I => \arses.counterZ0Z_1\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2582\,
            I => \arses.counterZ0Z_1\
        );

    \I__323\ : InMux
    port map (
            O => \N__2577\,
            I => \N__2571\
        );

    \I__322\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2568\
        );

    \I__321\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2563\
        );

    \I__320\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2563\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2571\,
            I => \arses.counterZ0Z_0\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2568\,
            I => \arses.counterZ0Z_0\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2563\,
            I => \arses.counterZ0Z_0\
        );

    \I__316\ : IoInMux
    port map (
            O => \N__2556\,
            I => \N__2553\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2553\,
            I => \N__2550\
        );

    \I__314\ : Odrv4
    port map (
            O => \N__2550\,
            I => lcol3_c
        );

    \I__313\ : CascadeMux
    port map (
            O => \N__2547\,
            I => \dig2.m13_am_cascade_\
        );

    \I__312\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2541\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2541\,
            I => \dig2.leds_17_i_0_ns_1_1\
        );

    \I__310\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2534\
        );

    \I__309\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2531\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2534\,
            I => \debounceup.counterZ0Z_3\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2531\,
            I => \debounceup.counterZ0Z_3\
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2526\,
            I => \debounceup.counter19_2_cascade_\
        );

    \I__305\ : InMux
    port map (
            O => \N__2523\,
            I => \N__2520\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2520\,
            I => \debounceup.counter_RNO_0_0_2\
        );

    \I__303\ : CascadeMux
    port map (
            O => \N__2517\,
            I => \debounceup.counter19_cascade_\
        );

    \I__302\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2510\
        );

    \I__301\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2507\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2510\,
            I => \debounceup.counterZ0Z_2\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2507\,
            I => \debounceup.counterZ0Z_2\
        );

    \I__298\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2492\
        );

    \I__297\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2492\
        );

    \I__296\ : InMux
    port map (
            O => \N__2500\,
            I => \N__2492\
        );

    \I__295\ : InMux
    port map (
            O => \N__2499\,
            I => \N__2489\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2492\,
            I => \N__2486\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2489\,
            I => \debounceup.counterZ0Z_4\
        );

    \I__292\ : Odrv4
    port map (
            O => \N__2486\,
            I => \debounceup.counterZ0Z_4\
        );

    \I__291\ : InMux
    port map (
            O => \N__2481\,
            I => \N__2476\
        );

    \I__290\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2471\
        );

    \I__289\ : InMux
    port map (
            O => \N__2479\,
            I => \N__2471\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2476\,
            I => \debounceup.counter19_2\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2471\,
            I => \debounceup.counter19_2\
        );

    \I__286\ : CascadeMux
    port map (
            O => \N__2466\,
            I => \dig2.m18_bm_cascade_\
        );

    \I__285\ : IoInMux
    port map (
            O => \N__2463\,
            I => \N__2460\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2460\,
            I => \N__2457\
        );

    \I__283\ : Span4Mux_s2_v
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__282\ : Span4Mux_v
    port map (
            O => \N__2454\,
            I => \N__2451\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__280\ : Span4Mux_v
    port map (
            O => \N__2448\,
            I => \N__2445\
        );

    \I__279\ : Odrv4
    port map (
            O => \N__2445\,
            I => leds_1_i_1
        );

    \I__278\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2438\
        );

    \I__277\ : InMux
    port map (
            O => \N__2441\,
            I => \N__2435\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2438\,
            I => \arses.counterZ0Z_7\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2435\,
            I => \arses.counterZ0Z_7\
        );

    \I__274\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2426\
        );

    \I__273\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2423\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2426\,
            I => \arses.counterZ0Z_6\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2423\,
            I => \arses.counterZ0Z_6\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__2418\,
            I => \N__2415\
        );

    \I__269\ : InMux
    port map (
            O => \N__2415\,
            I => \N__2411\
        );

    \I__268\ : InMux
    port map (
            O => \N__2414\,
            I => \N__2408\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2411\,
            I => \N__2405\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2408\,
            I => \arses.counterZ0Z_5\
        );

    \I__265\ : Odrv4
    port map (
            O => \N__2405\,
            I => \arses.counterZ0Z_5\
        );

    \I__264\ : InMux
    port map (
            O => \N__2400\,
            I => \N__2396\
        );

    \I__263\ : InMux
    port map (
            O => \N__2399\,
            I => \N__2393\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2396\,
            I => \arses.counterZ0Z_8\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2393\,
            I => \arses.counterZ0Z_8\
        );

    \I__260\ : InMux
    port map (
            O => \N__2388\,
            I => \N__2384\
        );

    \I__259\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2381\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2384\,
            I => \arses.counterZ0Z_3\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2381\,
            I => \arses.counterZ0Z_3\
        );

    \I__256\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2372\
        );

    \I__255\ : InMux
    port map (
            O => \N__2375\,
            I => \N__2369\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2372\,
            I => \arses.counterZ0Z_2\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2369\,
            I => \arses.counterZ0Z_2\
        );

    \I__252\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2360\
        );

    \I__251\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2357\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2360\,
            I => \arses.counterZ0Z_4\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2357\,
            I => \arses.counterZ0Z_4\
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2352\,
            I => \arses.un1_counterlto4_2_cascade_\
        );

    \I__247\ : InMux
    port map (
            O => \N__2349\,
            I => \N__2346\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2346\,
            I => \arses.un1_counterlto8_2\
        );

    \I__245\ : InMux
    port map (
            O => \N__2343\,
            I => \arses.un2_counter_cry_7\
        );

    \I__244\ : InMux
    port map (
            O => \N__2340\,
            I => \bfn_15_24_0_\
        );

    \I__243\ : InMux
    port map (
            O => \N__2337\,
            I => \arses.un2_counter_cry_9\
        );

    \I__242\ : InMux
    port map (
            O => \N__2334\,
            I => \arses.un2_counter_cry_10\
        );

    \I__241\ : InMux
    port map (
            O => \N__2331\,
            I => \arses.un2_counter_cry_11\
        );

    \I__240\ : InMux
    port map (
            O => \N__2328\,
            I => \arses.un2_counter_cry_12\
        );

    \I__239\ : InMux
    port map (
            O => \N__2325\,
            I => \arses.un2_counter_cry_13\
        );

    \I__238\ : IoInMux
    port map (
            O => \N__2322\,
            I => \N__2319\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2319\,
            I => \N__2316\
        );

    \I__236\ : IoSpan4Mux
    port map (
            O => \N__2316\,
            I => \N__2313\
        );

    \I__235\ : Span4Mux_s1_v
    port map (
            O => \N__2313\,
            I => \N__2310\
        );

    \I__234\ : Span4Mux_h
    port map (
            O => \N__2310\,
            I => \N__2307\
        );

    \I__233\ : Odrv4
    port map (
            O => \N__2307\,
            I => lcol4_c
        );

    \I__232\ : IoInMux
    port map (
            O => \N__2304\,
            I => \N__2301\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__2301\,
            I => \N__2298\
        );

    \I__230\ : IoSpan4Mux
    port map (
            O => \N__2298\,
            I => \N__2295\
        );

    \I__229\ : Odrv4
    port map (
            O => \N__2295\,
            I => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\
        );

    \I__228\ : InMux
    port map (
            O => \N__2292\,
            I => \debounceup.un3_counter_1_cry_2\
        );

    \I__227\ : InMux
    port map (
            O => \N__2289\,
            I => \debounceup.un3_counter_1_cry_3\
        );

    \I__226\ : InMux
    port map (
            O => \N__2286\,
            I => \arses.un2_counter_cry_1\
        );

    \I__225\ : InMux
    port map (
            O => \N__2283\,
            I => \arses.un2_counter_cry_2\
        );

    \I__224\ : InMux
    port map (
            O => \N__2280\,
            I => \arses.un2_counter_cry_3\
        );

    \I__223\ : InMux
    port map (
            O => \N__2277\,
            I => \arses.un2_counter_cry_4\
        );

    \I__222\ : InMux
    port map (
            O => \N__2274\,
            I => \arses.un2_counter_cry_5\
        );

    \I__221\ : InMux
    port map (
            O => \N__2271\,
            I => \arses.un2_counter_cry_6\
        );

    \I__220\ : IoInMux
    port map (
            O => \N__2268\,
            I => \N__2265\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2265\,
            I => \N__2262\
        );

    \I__218\ : IoSpan4Mux
    port map (
            O => \N__2262\,
            I => \N__2259\
        );

    \I__217\ : Span4Mux_s2_v
    port map (
            O => \N__2259\,
            I => \N__2256\
        );

    \I__216\ : Sp12to4
    port map (
            O => \N__2256\,
            I => \N__2253\
        );

    \I__215\ : Span12Mux_s10_v
    port map (
            O => \N__2253\,
            I => \N__2250\
        );

    \I__214\ : Span12Mux_v
    port map (
            O => \N__2250\,
            I => \N__2247\
        );

    \I__213\ : Span12Mux_h
    port map (
            O => \N__2247\,
            I => \N__2244\
        );

    \I__212\ : Odrv12
    port map (
            O => \N__2244\,
            I => \arse.divseven.io_0_D_IN_0\
        );

    \I__211\ : IoInMux
    port map (
            O => \N__2241\,
            I => \N__2238\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__2238\,
            I => \N__2235\
        );

    \I__209\ : Odrv4
    port map (
            O => \N__2235\,
            I => masterreset_c_i
        );

    \I__208\ : InMux
    port map (
            O => \N__2232\,
            I => \debounceup.un3_counter_1_cry_1\
        );

    \I__207\ : ClkMux
    port map (
            O => \N__2229\,
            I => \N__2226\
        );

    \I__206\ : GlobalMux
    port map (
            O => \N__2226\,
            I => \N__2223\
        );

    \I__205\ : gio2CtrlBuf
    port map (
            O => \N__2223\,
            I => \arse.un1_io_0_1_g\
        );

    \I__204\ : IoInMux
    port map (
            O => \N__2220\,
            I => \N__2217\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__2217\,
            I => \N__2214\
        );

    \I__202\ : IoSpan4Mux
    port map (
            O => \N__2214\,
            I => \N__2211\
        );

    \I__201\ : Span4Mux_s3_h
    port map (
            O => \N__2211\,
            I => \N__2208\
        );

    \I__200\ : Span4Mux_h
    port map (
            O => \N__2208\,
            I => \N__2205\
        );

    \I__199\ : Sp12to4
    port map (
            O => \N__2205\,
            I => \N__2202\
        );

    \I__198\ : Span12Mux_h
    port map (
            O => \N__2202\,
            I => \N__2199\
        );

    \I__197\ : Span12Mux_v
    port map (
            O => \N__2199\,
            I => \N__2196\
        );

    \I__196\ : Odrv12
    port map (
            O => \N__2196\,
            I => \top_pll_nrtthrth.PLLOUTCORE\
        );

    \INVarse.divseven.dout_0C\ : INV
    port map (
            O => \INVarse.divseven.dout_0C_net\,
            I => \N__5740\
        );

    \INVarse.apuresetoutregC\ : INV
    port map (
            O => \INVarse.apuresetoutregC_net\,
            I => \N__5747\
        );

    \INVarse.apusynclatchedC\ : INV
    port map (
            O => \INVarse.apusynclatchedC_net\,
            I => \N__2229\
        );

    \INVarse.diveight.dout_0C\ : INV
    port map (
            O => \INVarse.diveight.dout_0C_net\,
            I => \N__5749\
        );

    \INVarse.cpuclkresetC\ : INV
    port map (
            O => \INVarse.cpuclkresetC_net\,
            I => \N__5745\
        );

    \INVarse.cpuresetoutregC\ : INV
    port map (
            O => \INVarse.cpuresetoutregC_net\,
            I => \N__5751\
        );

    \INVarse.cpuresetcount_0C\ : INV
    port map (
            O => \INVarse.cpuresetcount_0C_net\,
            I => \N__5750\
        );

    \IN_MUX_bfv_27_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_27_10_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_24_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_17_0_\
        );

    \IN_MUX_bfv_20_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_17_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \arses.un2_counter_cry_8\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_29_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_29_7_0_\
        );

    \arses.clock_out_RNIR6ER_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2613\,
            GLOBALBUFFEROUTPUT => \N_111_g\
        );

    \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2220\,
            GLOBALBUFFEROUTPUT => \PLLOUTCORE_g\
        );

    \arse.divseven.io_0_RNIIG08\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2268\,
            GLOBALBUFFEROUTPUT => \arse.un1_io_0_1_g\
        );

    \masterreset_ibuf_RNIKP26_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2241\,
            GLOBALBUFFEROUTPUT => masterreset_c_i_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \masterreset_ibuf_RNIKP26_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => masterreset_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.un3_counter_1_cry_1_c_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3320\,
            in2 => \N__3347\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \debounceup.un3_counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_RNO_0_2_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2514\,
            in2 => \_gnd_net_\,
            in3 => \N__2232\,
            lcout => \debounceup.counter_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \debounceup.un3_counter_1_cry_1\,
            carryout => \debounceup.un3_counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_3_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2538\,
            in2 => \_gnd_net_\,
            in3 => \N__2292\,
            lcout => \debounceup.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \debounceup.un3_counter_1_cry_2\,
            carryout => \debounceup.un3_counter_1_cry_3\,
            clk => \N__4492\,
            ce => \N__4596\,
            sr => \_gnd_net_\
        );

    \debounceup.counter_4_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001000"
        )
    port map (
            in0 => \N__2499\,
            in1 => \N__2481\,
            in2 => \N__4652\,
            in3 => \N__2289\,
            lcout => \debounceup.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4492\,
            ce => \N__4596\,
            sr => \_gnd_net_\
        );

    \arses.un2_counter_cry_1_c_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2576\,
            in2 => \N__2598\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \arses.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_2_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2971\,
            in1 => \N__2376\,
            in2 => \_gnd_net_\,
            in3 => \N__2286\,
            lcout => \arses.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_1\,
            carryout => \arses.un2_counter_cry_2\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_3_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2963\,
            in1 => \N__2388\,
            in2 => \_gnd_net_\,
            in3 => \N__2283\,
            lcout => \arses.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_2\,
            carryout => \arses.un2_counter_cry_3\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_4_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2972\,
            in1 => \N__2364\,
            in2 => \_gnd_net_\,
            in3 => \N__2280\,
            lcout => \arses.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_3\,
            carryout => \arses.un2_counter_cry_4\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_5_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2964\,
            in1 => \N__2414\,
            in2 => \_gnd_net_\,
            in3 => \N__2277\,
            lcout => \arses.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_4\,
            carryout => \arses.un2_counter_cry_5\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_6_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2973\,
            in1 => \N__2430\,
            in2 => \_gnd_net_\,
            in3 => \N__2274\,
            lcout => \arses.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_5\,
            carryout => \arses.un2_counter_cry_6\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_7_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2965\,
            in1 => \N__2442\,
            in2 => \_gnd_net_\,
            in3 => \N__2271\,
            lcout => \arses.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_6\,
            carryout => \arses.un2_counter_cry_7\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_8_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2974\,
            in1 => \N__2400\,
            in2 => \_gnd_net_\,
            in3 => \N__2343\,
            lcout => \arses.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_7\,
            carryout => \arses.un2_counter_cry_8\,
            clk => \N__4506\,
            ce => 'H',
            sr => \N__4048\
        );

    \arses.counter_9_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2968\,
            in1 => \N__2667\,
            in2 => \_gnd_net_\,
            in3 => \N__2340\,
            lcout => \arses.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \arses.un2_counter_cry_9\,
            clk => \N__4509\,
            ce => 'H',
            sr => \N__4049\
        );

    \arses.counter_10_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2975\,
            in1 => \N__2682\,
            in2 => \_gnd_net_\,
            in3 => \N__2337\,
            lcout => \arses.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_9\,
            carryout => \arses.un2_counter_cry_10\,
            clk => \N__4509\,
            ce => 'H',
            sr => \N__4049\
        );

    \arses.counter_11_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2966\,
            in1 => \N__2694\,
            in2 => \_gnd_net_\,
            in3 => \N__2334\,
            lcout => \arses.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_10\,
            carryout => \arses.un2_counter_cry_11\,
            clk => \N__4509\,
            ce => 'H',
            sr => \N__4049\
        );

    \arses.counter_12_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2976\,
            in1 => \N__2628\,
            in2 => \_gnd_net_\,
            in3 => \N__2331\,
            lcout => \arses.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_11\,
            carryout => \arses.un2_counter_cry_12\,
            clk => \N__4509\,
            ce => 'H',
            sr => \N__4049\
        );

    \arses.counter_13_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2967\,
            in1 => \N__2643\,
            in2 => \_gnd_net_\,
            in3 => \N__2328\,
            lcout => \arses.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_12\,
            carryout => \arses.un2_counter_cry_13\,
            clk => \N__4509\,
            ce => 'H',
            sr => \N__4049\
        );

    \arses.counter_14_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2977\,
            in1 => \N__2655\,
            in2 => \_gnd_net_\,
            in3 => \N__2325\,
            lcout => \arses.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4509\,
            ce => 'H',
            sr => \N__4049\
        );

    \lcolreg_3_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__3581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3732\,
            lcout => lcol4_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4512\,
            ce => \N__4592\,
            sr => \_gnd_net_\
        );

    \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_RNI5J0P_2_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2537\,
            in2 => \_gnd_net_\,
            in3 => \N__2513\,
            lcout => \debounceup.counter19_2\,
            ltout => \debounceup.counter19_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_RNIADHU1_1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2500\,
            in1 => \N__3321\,
            in2 => \N__2526\,
            in3 => \N__3342\,
            lcout => \debounceup.counter19\,
            ltout => \debounceup.counter19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_2_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__2480\,
            in1 => \N__2523\,
            in2 => \N__2517\,
            in3 => \N__2502\,
            lcout => \debounceup.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4489\,
            ce => \N__4595\,
            sr => \_gnd_net_\
        );

    \debounceup.counter_0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__2501\,
            in1 => \N__2479\,
            in2 => \_gnd_net_\,
            in3 => \N__3343\,
            lcout => \debounceup.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4489\,
            ce => \N__4595\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m18_bm_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110001010"
        )
    port map (
            in0 => \N__4414\,
            in1 => \N__3572\,
            in2 => \N__4321\,
            in3 => \N__3095\,
            lcout => OPEN,
            ltout => \dig2.m18_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_1_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__4190\,
            in1 => \N__2733\,
            in2 => \N__2466\,
            in3 => \N__2544\,
            lcout => leds_1_i_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4489\,
            ce => \N__4595\,
            sr => \_gnd_net_\
        );

    \arses.counter_RNIA58_5_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2441\,
            in1 => \N__2429\,
            in2 => \N__2418\,
            in3 => \N__2399\,
            lcout => \arses.un1_counterlto8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI1L5_2_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2387\,
            in1 => \N__2375\,
            in2 => \_gnd_net_\,
            in3 => \N__2574\,
            lcout => OPEN,
            ltout => \arses.un1_counterlto4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOKH_1_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2363\,
            in1 => \N__2590\,
            in2 => \N__2352\,
            in3 => \N__2349\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI04C4_9_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2693\,
            in1 => \N__2681\,
            in2 => \N__2670\,
            in3 => \N__2666\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOS0A_14_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__2654\,
            in1 => \N__2642\,
            in2 => \N__2631\,
            in3 => \N__2627\,
            lcout => arses_counter8,
            ltout => \arses_counter8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_0_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4834\,
            in2 => \N__2616\,
            in3 => \N__2904\,
            lcout => \arses.clock_out_RNIR6ERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_1_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__2575\,
            in1 => \N__2970\,
            in2 => \_gnd_net_\,
            in3 => \N__2591\,
            lcout => \arses.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4503\,
            ce => 'H',
            sr => \N__4050\
        );

    \arses.counter_0_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2969\,
            in2 => \_gnd_net_\,
            in3 => \N__2577\,
            lcout => \arses.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4507\,
            ce => 'H',
            sr => \N__4052\
        );

    \lcolreg_2_LC_16_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3739\,
            in2 => \_gnd_net_\,
            in3 => \N__3571\,
            lcout => lcol3_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4511\,
            ce => \N__4591\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m13_am_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101001111010"
        )
    port map (
            in0 => \N__4412\,
            in1 => \N__3721\,
            in2 => \N__4311\,
            in3 => \N__3552\,
            lcout => OPEN,
            ltout => \dig2.m13_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_1_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__4181\,
            in1 => \N__4119\,
            in2 => \N__2547\,
            in3 => \N__2706\,
            lcout => \dig2.leds_17_i_0_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m18_am_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000100"
        )
    port map (
            in0 => \N__3553\,
            in1 => \N__4299\,
            in2 => \N__3738\,
            in3 => \N__4413\,
            lcout => \dig2.m18_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m77_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101100111111"
        )
    port map (
            in0 => \N__5615\,
            in1 => \N__3725\,
            in2 => \N__5315\,
            in3 => \N__3554\,
            lcout => \dig2.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_3_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__2700\,
            in1 => \N__4194\,
            in2 => \N__4110\,
            in3 => \N__2757\,
            lcout => leds_1_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4487\,
            ce => \N__4597\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m61_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101110100000"
        )
    port map (
            in0 => \N__5609\,
            in1 => \N__3659\,
            in2 => \N__5312\,
            in3 => \N__3476\,
            lcout => \dig2.i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m58_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110000100"
        )
    port map (
            in0 => \N__5610\,
            in1 => \N__3660\,
            in2 => \N__5311\,
            in3 => \N__3477\,
            lcout => \dig2.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m13_bm_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3478\,
            in1 => \N__4403\,
            in2 => \N__4295\,
            in3 => \N__3666\,
            lcout => \dig2.m13_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m41_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100101111111"
        )
    port map (
            in0 => \N__4384\,
            in1 => \N__3559\,
            in2 => \N__4322\,
            in3 => \N__3687\,
            lcout => \dig2.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m75_ns_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001010101"
        )
    port map (
            in0 => \N__2841\,
            in1 => \N__4996\,
            in2 => \N__3096\,
            in3 => \N__5614\,
            lcout => \dig2.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m54_am_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000010"
        )
    port map (
            in0 => \N__5611\,
            in1 => \N__3558\,
            in2 => \N__5313\,
            in3 => \N__3686\,
            lcout => \dig2.m54_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m69_am_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101001100111"
        )
    port map (
            in0 => \N__3560\,
            in1 => \N__5613\,
            in2 => \N__3720\,
            in3 => \N__5293\,
            lcout => \dig2.m69_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m69_bm_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001111000100"
        )
    port map (
            in0 => \N__5612\,
            in1 => \N__3561\,
            in2 => \N__5314\,
            in3 => \N__3691\,
            lcout => \dig2.m69_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_2_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010101"
        )
    port map (
            in0 => \N__2739\,
            in1 => \N__2835\,
            in2 => \N__2829\,
            in3 => \N__5689\,
            lcout => leds_1_i_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4490\,
            ce => \N__4598\,
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_0_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__3196\,
            in1 => \N__3182\,
            in2 => \_gnd_net_\,
            in3 => \N__3137\,
            lcout => \debounceconsolereset.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4490\,
            ce => \N__4598\,
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_1_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3161\,
            lcout => \debounceconsolereset.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4490\,
            ce => \N__4598\,
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_2_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__3240\,
            in1 => \N__3183\,
            in2 => \N__3201\,
            in3 => \N__3113\,
            lcout => \debounceconsolereset.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4490\,
            ce => \N__4598\,
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_3_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__2799\,
            in1 => \N__5690\,
            in2 => \N__2793\,
            in3 => \N__4997\,
            lcout => leds_1_i_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4490\,
            ce => \N__4598\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m39_ns_1_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110101"
        )
    port map (
            in0 => \N__4375\,
            in1 => \N__3658\,
            in2 => \N__4118\,
            in3 => \N__3475\,
            lcout => OPEN,
            ltout => \dig2.m39_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m39_ns_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000101"
        )
    port map (
            in0 => \N__4323\,
            in1 => \N__4114\,
            in2 => \N__2760\,
            in3 => \N__3087\,
            lcout => \dig2.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__2751\,
            in1 => \N__4995\,
            in2 => \N__5691\,
            in3 => \N__2745\,
            lcout => \dig2.leds_17_i_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m3_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3657\,
            in2 => \_gnd_net_\,
            in3 => \N__3474\,
            lcout => col_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \col_1_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__3091\,
            in1 => \N__3672\,
            in2 => \N__2903\,
            in3 => \N__3000\,
            lcout => \colZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_RNO_0_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2894\,
            in1 => \N__3112\,
            in2 => \N__4864\,
            in3 => \N__2987\,
            lcout => OPEN,
            ltout => \debounceconsolereset.out_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__3039\,
            in1 => \N__3024\,
            in2 => \N__3003\,
            in3 => \N__5387\,
            lcout => debouncedconsolereset,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__2986\,
            in1 => \N__4853\,
            in2 => \_gnd_net_\,
            in3 => \N__2893\,
            lcout => \clock_out_RNIR6ER\,
            ltout => \clock_out_RNIR6ER_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \col_0_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__2895\,
            in1 => \_gnd_net_\,
            in2 => \N__2994\,
            in3 => \N__3508\,
            lcout => \colZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__2991\,
            in1 => \N__4863\,
            in2 => \_gnd_net_\,
            in3 => \N__2899\,
            lcout => slowclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_1_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110010001"
        )
    port map (
            in0 => \N__5688\,
            in1 => \N__3048\,
            in2 => \N__2865\,
            in3 => \N__3057\,
            lcout => leds_1_i_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4491\,
            ce => \N__4601\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m75_ns_1_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110101"
        )
    port map (
            in0 => \N__5283\,
            in1 => \N__3692\,
            in2 => \N__4994\,
            in3 => \N__3557\,
            lcout => \dig2.m75_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_1_cry_1_c_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3136\,
            in2 => \N__3162\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_17_0_\,
            carryout => \debounceconsolereset.un3_counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNO_0_2_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3213\,
            in2 => \_gnd_net_\,
            in3 => \N__3234\,
            lcout => \debounceconsolereset.counter_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_1_cry_1\,
            carryout => \debounceconsolereset.un3_counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_3_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3225\,
            in2 => \_gnd_net_\,
            in3 => \N__3231\,
            lcout => \debounceconsolereset.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_1_cry_2\,
            carryout => \debounceconsolereset.un3_counter_1_cry_3\,
            clk => \N__4493\,
            ce => \N__4600\,
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_4_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001000"
        )
    port map (
            in0 => \N__3200\,
            in1 => \N__3181\,
            in2 => \N__3117\,
            in3 => \N__3228\,
            lcout => \debounceconsolereset.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4493\,
            ce => \N__4600\,
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNI7OV8_2_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3224\,
            in2 => \_gnd_net_\,
            in3 => \N__3212\,
            lcout => \debounceconsolereset.counter19_2\,
            ltout => \debounceconsolereset.counter19_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNIV9FM_1_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3180\,
            in1 => \N__3157\,
            in2 => \N__3141\,
            in3 => \N__3135\,
            lcout => \debounceconsolereset.counter19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m54_bm_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111010000"
        )
    port map (
            in0 => \N__5616\,
            in1 => \N__3488\,
            in2 => \N__5325\,
            in3 => \N__3086\,
            lcout => \dig2.m54_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_0_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__5282\,
            in1 => \N__4719\,
            in2 => \_gnd_net_\,
            in3 => \N__4758\,
            lcout => \delayConstantZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4488\,
            ce => 'H',
            sr => \N__4051\
        );

    \dig2.leds_cnst_3_1__leds_17_i_ns_1_1_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__4998\,
            in1 => \N__3294\,
            in2 => \N__5683\,
            in3 => \N__3288\,
            lcout => \dig2.leds_17_i_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_1_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3351\,
            in2 => \_gnd_net_\,
            in3 => \N__3313\,
            lcout => \debounceup.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4501\,
            ce => \N__4599\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m49_bm_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5586\,
            in1 => \N__3709\,
            in2 => \N__3586\,
            in3 => \N__5239\,
            lcout => \dig2.m49_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m33_am_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001010011011"
        )
    port map (
            in0 => \N__3579\,
            in1 => \N__4415\,
            in2 => \N__4303\,
            in3 => \N__3719\,
            lcout => \dig2.m33_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m49_am_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011100001010"
        )
    port map (
            in0 => \N__5587\,
            in1 => \N__3710\,
            in2 => \N__3587\,
            in3 => \N__5238\,
            lcout => \dig2.m49_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m33_bm_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010000111100"
        )
    port map (
            in0 => \N__4416\,
            in1 => \N__3737\,
            in2 => \N__3580\,
            in3 => \N__4294\,
            lcout => OPEN,
            ltout => \dig2.m33_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_2_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__4185\,
            in1 => \N__3282\,
            in2 => \N__3276\,
            in3 => \N__3252\,
            lcout => leds_1_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4496\,
            ce => \N__4603\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m22_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110000100"
        )
    port map (
            in0 => \N__4404\,
            in1 => \N__3736\,
            in2 => \N__4304\,
            in3 => \N__3556\,
            lcout => OPEN,
            ltout => \dig2.N_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__3246\,
            in1 => \N__4186\,
            in2 => \N__3255\,
            in3 => \N__4109\,
            lcout => \dig2.leds_17_i_0_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m25_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010001010"
        )
    port map (
            in0 => \N__3555\,
            in1 => \N__4405\,
            in2 => \N__3745\,
            in3 => \N__4285\,
            lcout => \dig2.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_0_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__3980\,
            in1 => \N__3956\,
            in2 => \_gnd_net_\,
            in3 => \N__3930\,
            lcout => \debouncedn.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4504\,
            ce => \N__4602\,
            sr => \_gnd_net_\
        );

    \lcolreg_0_LC_23_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3752\,
            in2 => \_gnd_net_\,
            in3 => \N__3591\,
            lcout => lcol1_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4513\,
            ce => \N__4594\,
            sr => \_gnd_net_\
        );

    \lcolreg_1_LC_23_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3753\,
            in2 => \_gnd_net_\,
            in3 => \N__3582\,
            lcout => lcol2_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4514\,
            ce => \N__4593\,
            sr => \_gnd_net_\
        );

    \debouncedn.counter_RNIVDIV_2_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3365\,
            in2 => \_gnd_net_\,
            in3 => \N__3386\,
            lcout => \debouncedn.counter19_2\,
            ltout => \debouncedn.counter19_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_RNIB0UE2_1_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3954\,
            in1 => \N__3933\,
            in2 => \N__3393\,
            in3 => \N__3903\,
            lcout => \debouncedn.counter19\,
            ltout => \debouncedn.counter19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_2_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__3957\,
            in1 => \N__3375\,
            in2 => \N__3390\,
            in3 => \N__3979\,
            lcout => \debouncedn.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4502\,
            ce => \N__4606\,
            sr => \_gnd_net_\
        );

    \debouncedn.un3_counter_1_cry_1_c_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3898\,
            in2 => \N__3932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_24_17_0_\,
            carryout => \debouncedn.un3_counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_RNO_0_2_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3387\,
            in2 => \_gnd_net_\,
            in3 => \N__3369\,
            lcout => \debouncedn.counter_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \debouncedn.un3_counter_1_cry_1\,
            carryout => \debouncedn.un3_counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_3_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3366\,
            in2 => \_gnd_net_\,
            in3 => \N__3354\,
            lcout => \debouncedn.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \debouncedn.un3_counter_1_cry_2\,
            carryout => \debouncedn.un3_counter_1_cry_3\,
            clk => \N__4505\,
            ce => \N__4605\,
            sr => \_gnd_net_\
        );

    \debouncedn.counter_4_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100000"
        )
    port map (
            in0 => \N__3955\,
            in1 => \N__3878\,
            in2 => \N__3984\,
            in3 => \N__3960\,
            lcout => \debouncedn.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4505\,
            ce => \N__4605\,
            sr => \_gnd_net_\
        );

    \debouncedn.counter_1_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3931\,
            in2 => \_gnd_net_\,
            in3 => \N__3902\,
            lcout => \debouncedn.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4508\,
            ce => \N__4604\,
            sr => \_gnd_net_\
        );

    \debouncedn.out_LC_26_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__3882\,
            in1 => \N__3864\,
            in2 => \N__4023\,
            in3 => \N__4614\,
            lcout => debounceddn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_26_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_0_c_LC_27_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4776\,
            in2 => \N__5326\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_27_10_0_\,
            carryout => \un1_delayConstant_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_1_LC_27_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4002\,
            in2 => \N__5571\,
            in3 => \N__3777\,
            lcout => \delayConstantZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_0\,
            carryout => \un1_delayConstant_cry_1\,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \delayConstant_2_LC_27_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4764\,
            in2 => \N__5649\,
            in3 => \N__3774\,
            lcout => \delayConstantZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_1\,
            carryout => \un1_delayConstant_cry_2\,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \delayConstant_3_LC_27_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4665\,
            in2 => \N__4971\,
            in3 => \N__3771\,
            lcout => \delayConstantZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_2\,
            carryout => \un1_delayConstant_cry_3\,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \delayConstant_4_LC_27_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3996\,
            in2 => \N__4374\,
            in3 => \N__4326\,
            lcout => \delayConstantZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_3\,
            carryout => \un1_delayConstant_cry_4\,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \delayConstant_5_LC_27_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3990\,
            in2 => \N__4259\,
            in3 => \N__4197\,
            lcout => \delayConstantZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_4\,
            carryout => \un1_delayConstant_cry_5\,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \delayConstant_6_LC_27_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4770\,
            in2 => \N__4171\,
            in3 => \N__4125\,
            lcout => \delayConstantZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_5\,
            carryout => \un1_delayConstant_cry_6\,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \delayConstant_7_LC_27_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__4706\,
            in1 => \N__4751\,
            in2 => \N__4089\,
            in3 => \N__4122\,
            lcout => \delayConstantZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4494\,
            ce => 'H',
            sr => \N__4053\
        );

    \olddn_LC_27_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4019\,
            lcout => \olddnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIEENH_LC_27_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4029\,
            in2 => \_gnd_net_\,
            in3 => \N__4018\,
            lcout => \olddn_RNIEENHZ0\,
            ltout => \olddn_RNIEENHZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_0_LC_27_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4005\,
            in3 => \N__4694\,
            lcout => \olddn_RNIM5BH1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_3_LC_28_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4748\,
            in1 => \_gnd_net_\,
            in2 => \N__4711\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNIM5BH1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_1_LC_28_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4702\,
            in2 => \_gnd_net_\,
            in3 => \N__4749\,
            lcout => \olddn_RNIM5BH1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oldup_RNI8NJV_LC_28_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__4852\,
            in1 => \N__4659\,
            in2 => \_gnd_net_\,
            in3 => \N__4541\,
            lcout => \delayConstant17_i\,
            ltout => \delayConstant17_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_0_c_RNO_LC_28_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \N__5327\,
            in1 => \_gnd_net_\,
            in2 => \N__4779\,
            in3 => \N__4745\,
            lcout => \un1_delayConstant_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_4_LC_28_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4750\,
            in1 => \_gnd_net_\,
            in2 => \N__4712\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNIM5BH1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_LC_28_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4695\,
            in2 => \_gnd_net_\,
            in3 => \N__4746\,
            lcout => \olddn_RNIM5BHZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_2_LC_28_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4747\,
            in1 => \_gnd_net_\,
            in2 => \N__4710\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNIM5BH1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oldup_LC_28_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4542\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \oldupZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.out_LC_28_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__4653\,
            in1 => \N__4632\,
            in2 => \N__4540\,
            in3 => \N__4613\,
            lcout => debouncedup,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_0_LC_29_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5172\,
            in2 => \N__5481\,
            in3 => \N__5480\,
            lcout => \arse.cpuresetcountZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_29_7_0_\,
            carryout => \arse.un1_cpuresetcount_1_cry_0\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_1_LC_29_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5138\,
            in2 => \_gnd_net_\,
            in3 => \N__4419\,
            lcout => \arse.cpuresetcountZ0Z_1\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_0\,
            carryout => \arse.un1_cpuresetcount_1_cry_1\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_2_LC_29_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5121\,
            in2 => \_gnd_net_\,
            in3 => \N__4914\,
            lcout => \arse.cpuresetcountZ0Z_2\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_1\,
            carryout => \arse.un1_cpuresetcount_1_cry_2\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_3_LC_29_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5055\,
            in2 => \_gnd_net_\,
            in3 => \N__4911\,
            lcout => \arse.cpuresetcountZ0Z_3\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_2\,
            carryout => \arse.un1_cpuresetcount_1_cry_3\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_4_LC_29_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5103\,
            in2 => \_gnd_net_\,
            in3 => \N__4908\,
            lcout => \arse.cpuresetcountZ0Z_4\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_3\,
            carryout => \arse.un1_cpuresetcount_1_cry_4\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_5_LC_29_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5156\,
            in2 => \_gnd_net_\,
            in3 => \N__4905\,
            lcout => \arse.cpuresetcountZ0Z_5\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_4\,
            carryout => \arse.un1_cpuresetcount_1_cry_5\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_6_LC_29_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5067\,
            in2 => \_gnd_net_\,
            in3 => \N__4902\,
            lcout => \arse.cpuresetcountZ0Z_6\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_5\,
            carryout => \arse.un1_cpuresetcount_1_cry_6\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \arse.cpuresetcount_7_LC_29_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5079\,
            in2 => \_gnd_net_\,
            in3 => \N__4899\,
            lcout => \arse.cpuresetcountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5028\
        );

    \debounceconsolereset.out_RNI1B6C_LC_29_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => debouncedconsolereset_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_LC_30_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4892\,
            in2 => \_gnd_net_\,
            in3 => \N__5085\,
            lcout => \arse.cpuresetoutregZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuresetoutregC_net\,
            ce => 'H',
            sr => \N__5027\
        );

    \arse.cpuclkreset_RNO_1_LC_30_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5119\,
            in1 => \N__5170\,
            in2 => \N__5157\,
            in3 => \N__5134\,
            lcout => OPEN,
            ltout => \arse.m8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuclkreset_RNO_0_LC_30_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5469\,
            in1 => \N__5101\,
            in2 => \N__5175\,
            in3 => \N__5042\,
            lcout => \arse.cpuclkreset_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_1_LC_30_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5171\,
            in1 => \N__5155\,
            in2 => \N__5139\,
            in3 => \N__5120\,
            lcout => OPEN,
            ltout => \arse.m12_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_0_LC_30_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5043\,
            in1 => \N__5470\,
            in2 => \N__5106\,
            in3 => \N__5102\,
            lcout => \arse.cpuresetoutreg_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_RNIFLN61_7_LC_30_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5078\,
            in1 => \N__5066\,
            in2 => \_gnd_net_\,
            in3 => \N__5054\,
            lcout => \arse.m4_e_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuclkreset_LC_30_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5034\,
            in2 => \_gnd_net_\,
            in3 => \N__5516\,
            lcout => arse_cpuclkreset,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuclkresetC_net\,
            ce => 'H',
            sr => \N__5026\
        );

    \arse.diveight.dout_0_LC_31_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5206\,
            in2 => \_gnd_net_\,
            in3 => \N__5520\,
            lcout => \arse.diveight.doutZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.diveight.dout_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_RNI7BAS_1_LC_31_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5368\,
            in2 => \_gnd_net_\,
            in3 => \N__5352\,
            lcout => OPEN,
            ltout => \arse_diveight_N_123_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_2_LC_31_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__4990\,
            in1 => \N__5207\,
            in2 => \N__4917\,
            in3 => \N__5514\,
            lcout => arse_diveight_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_1_LC_31_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__5513\,
            in1 => \N__5369\,
            in2 => \N__5684\,
            in3 => \N__5353\,
            lcout => arse_diveight_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5746\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_RNO_1_LC_31_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5512\,
            lcout => \arse.diveight.cpuclkreset_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_0_LC_31_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__5588\,
            in1 => \N__5355\,
            in2 => \_gnd_net_\,
            in3 => \N__5515\,
            lcout => arse_diveight_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.apusynclatched_LC_32_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__5487\,
            in1 => \N__5453\,
            in2 => \_gnd_net_\,
            in3 => \N__5424\,
            lcout => \arse.apusynclatchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.apusynclatchedC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.io_0_RNO_0_LC_32_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \arse.diveight.dout_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.io_0_RNO_LC_32_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5190\,
            lcout => \arse.diveight.dout_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.apuresetoutreg_LC_32_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5420\,
            lcout => \arse.apuresetoutregZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.apuresetoutregC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_1_LC_32_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__5370\,
            in1 => \N__5354\,
            in2 => \N__5334\,
            in3 => \N__5208\,
            lcout => \arse.diveight.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5743\,
            ce => 'H',
            sr => \N__5184\
        );

    \arse.divseven.counter_2_LC_32_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__5811\,
            in1 => \N__5799\,
            in2 => \_gnd_net_\,
            in3 => \N__5768\,
            lcout => \arse.divseven.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_1_LC_32_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5810\,
            in2 => \_gnd_net_\,
            in3 => \N__5798\,
            lcout => \arse.divseven.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_0_LC_32_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5797\,
            lcout => \arse.divseven.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_0_LC_32_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5767\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \arse.divseven.doutZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.divseven.dout_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.io_0_RNO_0_LC_32_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5787\,
            in3 => \_gnd_net_\,
            lcout => \arse.divseven.dout_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_1_LC_32_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5772\,
            lcout => \arse.divseven.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.io_0_RNO_LC_32_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5703\,
            lcout => \arse.divseven.dout_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
