// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 11 2024 23:52:07

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    masterreset,
    led4,
    lcol3,
    led5,
    lcol2,
    led6,
    led2,
    lcol1,
    deldn,
    cpuclk,
    apureset,
    led7,
    led3,
    lcol4,
    delup,
    cpureset,
    apusync,
    PACKAGEPIN,
    led8,
    led1,
    consolereset,
    apuclk);

    input masterreset;
    output led4;
    output lcol3;
    output led5;
    output lcol2;
    output led6;
    output led2;
    output lcol1;
    input deldn;
    output cpuclk;
    output apureset;
    output led7;
    output led3;
    output lcol4;
    input delup;
    output cpureset;
    input apusync;
    input PACKAGEPIN;
    output led8;
    output led1;
    input consolereset;
    output apuclk;

    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6465;
    wire N__6464;
    wire N__6463;
    wire N__6456;
    wire N__6455;
    wire N__6454;
    wire N__6447;
    wire N__6446;
    wire N__6445;
    wire N__6438;
    wire N__6437;
    wire N__6436;
    wire N__6429;
    wire N__6428;
    wire N__6427;
    wire N__6420;
    wire N__6419;
    wire N__6418;
    wire N__6411;
    wire N__6410;
    wire N__6409;
    wire N__6402;
    wire N__6401;
    wire N__6400;
    wire N__6393;
    wire N__6392;
    wire N__6391;
    wire N__6384;
    wire N__6383;
    wire N__6382;
    wire N__6375;
    wire N__6374;
    wire N__6373;
    wire N__6366;
    wire N__6365;
    wire N__6364;
    wire N__6357;
    wire N__6356;
    wire N__6355;
    wire N__6348;
    wire N__6347;
    wire N__6346;
    wire N__6339;
    wire N__6338;
    wire N__6337;
    wire N__6330;
    wire N__6329;
    wire N__6328;
    wire N__6321;
    wire N__6320;
    wire N__6319;
    wire N__6312;
    wire N__6311;
    wire N__6310;
    wire N__6303;
    wire N__6302;
    wire N__6301;
    wire N__6294;
    wire N__6293;
    wire N__6292;
    wire N__6285;
    wire N__6284;
    wire N__6283;
    wire N__6266;
    wire N__6265;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6257;
    wire N__6256;
    wire N__6255;
    wire N__6252;
    wire N__6245;
    wire N__6240;
    wire N__6233;
    wire N__6232;
    wire N__6231;
    wire N__6230;
    wire N__6229;
    wire N__6226;
    wire N__6225;
    wire N__6222;
    wire N__6211;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6190;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6175;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6157;
    wire N__6154;
    wire N__6153;
    wire N__6148;
    wire N__6145;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6107;
    wire N__6104;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6066;
    wire N__6065;
    wire N__6062;
    wire N__6055;
    wire N__6050;
    wire N__6049;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6041;
    wire N__6040;
    wire N__6039;
    wire N__6036;
    wire N__6031;
    wire N__6024;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6010;
    wire N__6009;
    wire N__6006;
    wire N__6001;
    wire N__5996;
    wire N__5993;
    wire N__5992;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5939;
    wire N__5934;
    wire N__5927;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5915;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5911;
    wire N__5910;
    wire N__5909;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5902;
    wire N__5901;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5841;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5785;
    wire N__5784;
    wire N__5781;
    wire N__5780;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5765;
    wire N__5760;
    wire N__5759;
    wire N__5756;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5738;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5730;
    wire N__5729;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5712;
    wire N__5709;
    wire N__5708;
    wire N__5705;
    wire N__5698;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5683;
    wire N__5680;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5662;
    wire N__5661;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5548;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5516;
    wire N__5513;
    wire N__5512;
    wire N__5509;
    wire N__5508;
    wire N__5507;
    wire N__5506;
    wire N__5503;
    wire N__5502;
    wire N__5497;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5490;
    wire N__5489;
    wire N__5486;
    wire N__5481;
    wire N__5478;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5450;
    wire N__5447;
    wire N__5442;
    wire N__5437;
    wire N__5432;
    wire N__5423;
    wire N__5420;
    wire N__5419;
    wire N__5418;
    wire N__5417;
    wire N__5416;
    wire N__5415;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5407;
    wire N__5406;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5386;
    wire N__5385;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5371;
    wire N__5366;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5344;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5322;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5308;
    wire N__5307;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5285;
    wire N__5282;
    wire N__5281;
    wire N__5280;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5212;
    wire N__5211;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5190;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5180;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5162;
    wire N__5159;
    wire N__5158;
    wire N__5155;
    wire N__5154;
    wire N__5153;
    wire N__5152;
    wire N__5151;
    wire N__5148;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5112;
    wire N__5107;
    wire N__5102;
    wire N__5093;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5087;
    wire N__5084;
    wire N__5083;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5032;
    wire N__5021;
    wire N__5020;
    wire N__5017;
    wire N__5016;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5004;
    wire N__4997;
    wire N__4996;
    wire N__4995;
    wire N__4994;
    wire N__4993;
    wire N__4990;
    wire N__4983;
    wire N__4980;
    wire N__4973;
    wire N__4972;
    wire N__4969;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4841;
    wire N__4840;
    wire N__4839;
    wire N__4838;
    wire N__4837;
    wire N__4836;
    wire N__4835;
    wire N__4834;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4786;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4782;
    wire N__4781;
    wire N__4780;
    wire N__4779;
    wire N__4778;
    wire N__4777;
    wire N__4776;
    wire N__4775;
    wire N__4774;
    wire N__4773;
    wire N__4772;
    wire N__4771;
    wire N__4770;
    wire N__4769;
    wire N__4768;
    wire N__4767;
    wire N__4766;
    wire N__4765;
    wire N__4764;
    wire N__4763;
    wire N__4762;
    wire N__4761;
    wire N__4760;
    wire N__4757;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4682;
    wire N__4681;
    wire N__4680;
    wire N__4679;
    wire N__4678;
    wire N__4675;
    wire N__4670;
    wire N__4667;
    wire N__4666;
    wire N__4665;
    wire N__4664;
    wire N__4663;
    wire N__4662;
    wire N__4661;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4640;
    wire N__4639;
    wire N__4638;
    wire N__4637;
    wire N__4634;
    wire N__4633;
    wire N__4630;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4619;
    wire N__4618;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4606;
    wire N__4601;
    wire N__4596;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4588;
    wire N__4587;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4572;
    wire N__4569;
    wire N__4564;
    wire N__4557;
    wire N__4554;
    wire N__4549;
    wire N__4544;
    wire N__4539;
    wire N__4530;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4489;
    wire N__4488;
    wire N__4485;
    wire N__4480;
    wire N__4477;
    wire N__4476;
    wire N__4475;
    wire N__4474;
    wire N__4473;
    wire N__4472;
    wire N__4471;
    wire N__4470;
    wire N__4467;
    wire N__4466;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4460;
    wire N__4455;
    wire N__4454;
    wire N__4453;
    wire N__4452;
    wire N__4451;
    wire N__4450;
    wire N__4449;
    wire N__4448;
    wire N__4447;
    wire N__4446;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4440;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4421;
    wire N__4416;
    wire N__4411;
    wire N__4406;
    wire N__4401;
    wire N__4394;
    wire N__4389;
    wire N__4382;
    wire N__4377;
    wire N__4352;
    wire N__4351;
    wire N__4350;
    wire N__4349;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4337;
    wire N__4336;
    wire N__4335;
    wire N__4334;
    wire N__4333;
    wire N__4332;
    wire N__4331;
    wire N__4330;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4322;
    wire N__4319;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4311;
    wire N__4310;
    wire N__4309;
    wire N__4308;
    wire N__4307;
    wire N__4306;
    wire N__4305;
    wire N__4304;
    wire N__4301;
    wire N__4296;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4271;
    wire N__4266;
    wire N__4259;
    wire N__4254;
    wire N__4247;
    wire N__4240;
    wire N__4217;
    wire N__4216;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4212;
    wire N__4209;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4201;
    wire N__4198;
    wire N__4197;
    wire N__4196;
    wire N__4195;
    wire N__4192;
    wire N__4187;
    wire N__4184;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4141;
    wire N__4132;
    wire N__4129;
    wire N__4118;
    wire N__4115;
    wire N__4114;
    wire N__4113;
    wire N__4112;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4051;
    wire N__4050;
    wire N__4049;
    wire N__4048;
    wire N__4047;
    wire N__4046;
    wire N__4041;
    wire N__4040;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4033;
    wire N__4028;
    wire N__4023;
    wire N__4020;
    wire N__4015;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__3999;
    wire N__3992;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3913;
    wire N__3912;
    wire N__3911;
    wire N__3908;
    wire N__3907;
    wire N__3906;
    wire N__3905;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3891;
    wire N__3884;
    wire N__3875;
    wire N__3874;
    wire N__3873;
    wire N__3872;
    wire N__3871;
    wire N__3870;
    wire N__3869;
    wire N__3868;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3854;
    wire N__3845;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3820;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3812;
    wire N__3811;
    wire N__3808;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3788;
    wire N__3787;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3691;
    wire N__3690;
    wire N__3687;
    wire N__3682;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3585;
    wire N__3584;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3560;
    wire N__3559;
    wire N__3554;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3505;
    wire N__3504;
    wire N__3501;
    wire N__3496;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3418;
    wire N__3417;
    wire N__3416;
    wire N__3415;
    wire N__3414;
    wire N__3413;
    wire N__3412;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3398;
    wire N__3397;
    wire N__3390;
    wire N__3381;
    wire N__3374;
    wire N__3367;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3332;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3293;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3278;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3266;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3254;
    wire N__3253;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3230;
    wire N__3227;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3215;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3203;
    wire N__3200;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3188;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3176;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3164;
    wire N__3161;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3149;
    wire N__3146;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3134;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3112;
    wire N__3111;
    wire N__3108;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3049;
    wire N__3048;
    wire N__3047;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3029;
    wire N__3028;
    wire N__3027;
    wire N__3026;
    wire N__3021;
    wire N__3016;
    wire N__3011;
    wire N__3010;
    wire N__3009;
    wire N__3006;
    wire N__3001;
    wire N__2996;
    wire N__2993;
    wire N__2992;
    wire N__2989;
    wire N__2988;
    wire N__2985;
    wire N__2984;
    wire N__2981;
    wire N__2974;
    wire N__2969;
    wire N__2966;
    wire N__2965;
    wire N__2962;
    wire N__2961;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2949;
    wire N__2942;
    wire N__2941;
    wire N__2940;
    wire N__2935;
    wire N__2932;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2869;
    wire N__2868;
    wire N__2865;
    wire N__2860;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2842;
    wire N__2841;
    wire N__2838;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2826;
    wire N__2823;
    wire N__2816;
    wire N__2815;
    wire N__2812;
    wire N__2811;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2799;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2782;
    wire N__2781;
    wire N__2780;
    wire N__2777;
    wire N__2772;
    wire N__2769;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2734;
    wire N__2733;
    wire N__2728;
    wire N__2725;
    wire N__2720;
    wire N__2719;
    wire N__2716;
    wire N__2715;
    wire N__2714;
    wire N__2711;
    wire N__2704;
    wire N__2701;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2686;
    wire N__2685;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2673;
    wire N__2670;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2653;
    wire N__2652;
    wire N__2651;
    wire N__2648;
    wire N__2643;
    wire N__2640;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2626;
    wire N__2623;
    wire N__2622;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2610;
    wire N__2603;
    wire N__2602;
    wire N__2601;
    wire N__2600;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2573;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2494;
    wire N__2493;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2477;
    wire N__2476;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2456;
    wire N__2453;
    wire N__2450;
    wire N__2447;
    wire N__2444;
    wire N__2441;
    wire N__2438;
    wire N__2435;
    wire N__2432;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2417;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire \arse.un1_io_0_1_g ;
    wire \top_pll_nrtthrth.PLLOUTCORE ;
    wire GNDG0;
    wire \arse.divseven.io_0_D_IN_0 ;
    wire VCCG0;
    wire masterreset_c_i;
    wire bfn_15_15_0_;
    wire \debouncedn.un3_counter_cry_1 ;
    wire \debouncedn.un3_counter_cry_2 ;
    wire \debouncedn.un3_counter_cry_3 ;
    wire GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO;
    wire \debouncedn.counter18_0_2_cascade_ ;
    wire \debouncedn.counterZ0Z_1 ;
    wire \debouncedn.counterZ0Z_4 ;
    wire \debouncedn.counter_RNIBTPA2Z0Z_4_cascade_ ;
    wire \debouncedn.counterZ0Z_0 ;
    wire \debounceconsolereset.counter18_0_2_cascade_ ;
    wire \debouncedn.un3_counter_cry_2_THRU_CO ;
    wire \debouncedn.counterZ0Z_3 ;
    wire \debouncedn.un3_counter_cry_1_THRU_CO ;
    wire \debouncedn.counter_RNIBTPA2Z0Z_4 ;
    wire \debouncedn.counterZ0Z_2 ;
    wire consolereset_c;
    wire \debounceconsolereset.out_cnv_2 ;
    wire lcol3_c;
    wire lcol4_c;
    wire bfn_17_14_0_;
    wire \debounceup.un3_counter_cry_1 ;
    wire \debounceup.un3_counter_cry_2 ;
    wire \debounceup.un3_counter_cry_3 ;
    wire \debounceup.un3_counter_cry_2_THRU_CO ;
    wire \debounceup.un3_counter_cry_1_THRU_CO ;
    wire \debounceconsolereset.counterZ0Z_1 ;
    wire \debounceconsolereset.counterZ0Z_0 ;
    wire bfn_17_15_0_;
    wire \debounceconsolereset.un3_counter_cry_1 ;
    wire \debounceconsolereset.un3_counter_cry_2 ;
    wire \debounceconsolereset.un3_counter_cry_3 ;
    wire \debounceconsolereset.counterZ0Z_4 ;
    wire clock_out_RNIR6ER_0_cascade_;
    wire \debounceconsolereset.un3_counter_cry_2_THRU_CO ;
    wire \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_ ;
    wire \debounceconsolereset.counterZ0Z_3 ;
    wire \debounceconsolereset.counter_RNINST81Z0Z_4 ;
    wire \debounceconsolereset.un3_counter_cry_1_THRU_CO ;
    wire \debounceconsolereset.counterZ0Z_2 ;
    wire bfn_17_16_0_;
    wire \arses.un2_counter_cry_1 ;
    wire \arses.un2_counter_cry_2 ;
    wire \arses.un2_counter_cry_3 ;
    wire \arses.un2_counter_cry_4 ;
    wire \arses.un2_counter_cry_5 ;
    wire \arses.un2_counter_cry_6 ;
    wire \arses.un2_counter_cry_7 ;
    wire \arses.un2_counter_cry_8 ;
    wire bfn_17_17_0_;
    wire \arses.un2_counter_cry_9 ;
    wire \arses.un2_counter_cry_10 ;
    wire \arses.un2_counter_cry_11 ;
    wire \arses.un2_counter_cry_12 ;
    wire \arses.un2_counter_cry_13 ;
    wire leds_1_i_0_3;
    wire \debounceup.counter_RNI45V02Z0Z_4_cascade_ ;
    wire \debounceup.counterZ0Z_3 ;
    wire \debounceup.counterZ0Z_2 ;
    wire \debounceup.counterZ0Z_4 ;
    wire \debounceup.counter18_0_2_cascade_ ;
    wire \debounceup.counterZ0Z_0 ;
    wire \debounceup.counter_RNI45V02Z0Z_4 ;
    wire \debounceup.counterZ0Z_1 ;
    wire leds_1_i_0_2;
    wire \arses.counterZ0Z_7 ;
    wire \arses.counterZ0Z_6 ;
    wire \arses.counterZ0Z_8 ;
    wire \arses.counterZ0Z_5 ;
    wire \arses.counterZ0Z_4 ;
    wire \arses.counterZ0Z_1 ;
    wire \arses.un1_counterlto8_2_cascade_ ;
    wire \arses.counterZ0Z_11 ;
    wire \arses.counterZ0Z_10 ;
    wire \arses.un1_counterlt11_cascade_ ;
    wire \arses.counterZ0Z_9 ;
    wire \arses.counterZ0Z_14 ;
    wire \arses.counterZ0Z_13 ;
    wire \arses.un1_counterlt13_0_cascade_ ;
    wire \arses.counterZ0Z_12 ;
    wire \arses.counter8_cascade_ ;
    wire \arses.counterZ0Z_3 ;
    wire \arses.counterZ0Z_2 ;
    wire \arses.un1_counterlto4_2 ;
    wire \arses.counterZ0Z_0 ;
    wire \dig1.N_78 ;
    wire \dig1.N_72 ;
    wire \debouncedn.out_cnv_2 ;
    wire deldn_c;
    wire \dig1.N_58_cascade_ ;
    wire \dig1.leds_17_i_ns_1_2 ;
    wire \dig1.N_61 ;
    wire \dig1.m68_bm ;
    wire \dig1.m68_am ;
    wire \arses.counter8 ;
    wire lcol2_c;
    wire masterreset_c;
    wire delayConstant16_i_cascade_;
    wire oldupZ0;
    wire debounceddn;
    wire olddnZ0;
    wire \dig1.m77_am ;
    wire \debounceup.out_cnv_2 ;
    wire delup_c;
    wire debouncedup;
    wire \dig1.m77_bm ;
    wire leds_1_i_1;
    wire lcol1_c;
    wire \dig1.N_39 ;
    wire leds_1_i_3;
    wire \dig1.N_15_cascade_ ;
    wire \dig1.N_18 ;
    wire slowclk;
    wire clock_out_RNIR6ER;
    wire \dig1.N_17 ;
    wire \dig1.m32_bm ;
    wire \dig1.m32_am ;
    wire leds_1_i_2;
    wire un1_delayConstant_cry_0_c_RNOZ0;
    wire bfn_21_12_0_;
    wire olddn_RNIM5BH1Z0Z_1;
    wire un1_delayConstant_cry_0;
    wire olddn_RNIM5BHZ0Z1;
    wire un1_delayConstant_cry_1;
    wire olddn_RNIM5BH1Z0Z_2;
    wire un1_delayConstant_cry_2;
    wire olddn_RNIM5BH1Z0Z_3;
    wire un1_delayConstant_cry_3;
    wire olddn_RNIM5BH1Z0Z_0;
    wire un1_delayConstant_cry_4;
    wire olddn_RNIM5BH1Z0Z_4;
    wire un1_delayConstant_cry_5;
    wire delayConstant16_i;
    wire olddn_RNIEENHZ0;
    wire un1_delayConstant_cry_6;
    wire \dig1.m41_bm ;
    wire \dig1.m41_am_cascade_ ;
    wire \dig1.N_44 ;
    wire \dig1.m10_ns_1_cascade_ ;
    wire \dig1.N_11_0 ;
    wire delayConstantZ0Z_6;
    wire \dig1.N_25 ;
    wire \dig1.N_22_cascade_ ;
    wire \dig1.leds_17_i_0_ns_1_2 ;
    wire un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2;
    wire un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92;
    wire masterreset_c_i_g;
    wire leds_1_i_0_1;
    wire PACKAGEPIN_0_c_g;
    wire clock_out_RNIR6ER_0;
    wire \dig1.N_52_cascade_ ;
    wire \dig1.N_54 ;
    wire \dig1.N_55 ;
    wire colZ0Z_0;
    wire colZ0Z_1;
    wire delayConstantZ0Z_2;
    wire \dig1.m47_ns_1_cascade_ ;
    wire col_1_1;
    wire \dig1.N_49 ;
    wire CONSTANT_ONE_NET;
    wire bfn_27_8_0_;
    wire \arse.un1_cpuresetcount_1_cry_0 ;
    wire \arse.un1_cpuresetcount_1_cry_1 ;
    wire \arse.un1_cpuresetcount_1_cry_2 ;
    wire \arse.un1_cpuresetcount_1_cry_3 ;
    wire \arse.un1_cpuresetcount_1_cry_4 ;
    wire \arse.un1_cpuresetcount_1_cry_5 ;
    wire \arse.un1_cpuresetcount_1_cry_6 ;
    wire \INVarse.cpuresetcount_0C_net ;
    wire delayConstantZ0Z_1;
    wire delayConstantZ0Z_5;
    wire \arse.g0_i_a3_4 ;
    wire \arse.cpuresetcountZ0Z_5 ;
    wire \arse.doingseven3_6_cascade_ ;
    wire \arse.cpuresetcountZ0Z_1 ;
    wire \arse.doingseven3_1 ;
    wire \arse.doingseven3_6 ;
    wire \arse.doingseven3_1_cascade_ ;
    wire delayConstant_fastZ0Z_6;
    wire delayConstant_fastZ0Z_2;
    wire \arse.cpuresetcountZ0Z_6 ;
    wire \arse.cpuresetcountZ0Z_2 ;
    wire delayConstantZ0Z_7;
    wire delayConstantZ0Z_3;
    wire \arse.cpuresetcountZ0Z_7 ;
    wire \arse.cpuresetcountZ0Z_3 ;
    wire delayConstantZ0Z_4;
    wire delayConstantZ0Z_0;
    wire \arse.cpuresetcountZ0Z_0 ;
    wire \arse.cpuresetcountZ0Z_4 ;
    wire \arse.g0_3 ;
    wire \arse.g0_2_cascade_ ;
    wire \arse.g0_4 ;
    wire \arse.N_6 ;
    wire \arse.g0_1 ;
    wire \arse.g0_7_cascade_ ;
    wire \arse.cpuresetoutreg_1_sqmuxa_cascade_ ;
    wire \arse.cpuresetoutregZ0 ;
    wire \INVarse.cpuresetoutregC_net ;
    wire \arse.doingseven4 ;
    wire \INVarse.cpuclkresetC_net ;
    wire \arse.doingseven3 ;
    wire \INVarse.doingsevenC_net ;
    wire debouncedconsolereset_i;
    wire \arse.doingsevenZ0 ;
    wire \arse.diveight.doutZ1Z_0 ;
    wire \INVarse.diveight.dout_0C_net ;
    wire \arse.divseven.un1_counter_i_0_0 ;
    wire \arse.divseven.counterZ0Z_0 ;
    wire \arse.divseven.sevenZ0 ;
    wire apusync_c;
    wire \arse.apusynclatchedZ0 ;
    wire \INVarse.apusynclatchedC_net ;
    wire debouncedconsolereset;
    wire \arse.apuresetoutregZ0 ;
    wire \INVarse.apuresetoutregC_net ;
    wire \arse.diveight.counterZ0Z_0 ;
    wire \arse.cpuclkresetZ0 ;
    wire \arse.diveight.counterZ0Z_1 ;
    wire \arse.diveight.counterZ0Z_2 ;
    wire \arse.diveight.doutZ0Z_1 ;
    wire \arse.divseven.N_46_0 ;
    wire \arse.divseven.counterZ0Z_1 ;
    wire \arse.divseven.doutZ0Z_1 ;
    wire PLLOUTCORE_g;
    wire \arse.divseven.counterZ0Z_2 ;
    wire \arse.divseven.doutZ0Z_0 ;
    wire \INVarse.divseven.dout_0C_net ;
    wire \arse.divseven.un1_dout_2_sqmuxa_0_i ;
    wire _gnd_net_;

    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .TEST_MODE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FILTER_RANGE=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_RELATIVE=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVR=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVQ=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVF=7'b0011111;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \top_pll_nrtthrth.top_pll_nrtthrth_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\top_pll_nrtthrth.PLLOUTCORE ),
            .REFERENCECLK(N__2510),
            .RESETB(N__3602),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF PACKAGEPIN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6474),
            .GLOBALBUFFEROUTPUT(PACKAGEPIN_0_c_g));
    IO_PAD PACKAGEPIN_ibuf_gb_io_iopad (
            .OE(N__6476),
            .DIN(N__6475),
            .DOUT(N__6474),
            .PACKAGEPIN(PACKAGEPIN));
    defparam PACKAGEPIN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam PACKAGEPIN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO PACKAGEPIN_ibuf_gb_io_preio (
            .PADOEN(N__6476),
            .PADOUT(N__6475),
            .PADIN(N__6474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD masterreset_ibuf_iopad (
            .OE(N__6465),
            .DIN(N__6464),
            .DOUT(N__6463),
            .PACKAGEPIN(masterreset));
    defparam masterreset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam masterreset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO masterreset_ibuf_preio (
            .PADOEN(N__6465),
            .PADOUT(N__6464),
            .PADIN(N__6463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(masterreset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led3_obuf_iopad (
            .OE(N__6456),
            .DIN(N__6455),
            .DOUT(N__6454),
            .PACKAGEPIN(led3));
    defparam led3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led3_obuf_preio (
            .PADOEN(N__6456),
            .PADOUT(N__6455),
            .PADIN(N__6454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2927),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.divseven.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.divseven.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.divseven.io_0_iopad  (
            .OE(N__6447),
            .DIN(N__6446),
            .DOUT(N__6445),
            .PACKAGEPIN(apuclk));
    defparam \arse.divseven.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.divseven.io_0_preio  (
            .PADOEN(N__6447),
            .PADOUT(N__6446),
            .PADIN(N__6445),
            .CLOCKENABLE(),
            .DOUT1(N__5926),
            .OUTPUTENABLE(N__4973),
            .DIN0(\arse.divseven.io_0_D_IN_0 ),
            .DOUT0(N__5834),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5909));
    defparam \arse.io_1_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.io_1_iopad .PULLUP=1'b0;
    IO_PAD \arse.io_1_iopad  (
            .OE(N__6438),
            .DIN(N__6437),
            .DOUT(N__6436),
            .PACKAGEPIN(cpureset));
    defparam \arse.io_1_preio .PIN_TYPE=6'b010101;
    PRE_IO \arse.io_1_preio  (
            .PADOEN(N__6438),
            .PADOUT(N__6437),
            .PADIN(N__6436),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5579),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5915));
    IO_PAD lcol3_obuf_iopad (
            .OE(N__6429),
            .DIN(N__6428),
            .DOUT(N__6427),
            .PACKAGEPIN(lcol3));
    defparam lcol3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol3_obuf_preio (
            .PADOEN(N__6429),
            .PADOUT(N__6428),
            .PADIN(N__6427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2555),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD deldn_ibuf_iopad (
            .OE(N__6420),
            .DIN(N__6419),
            .DOUT(N__6418),
            .PACKAGEPIN(deldn));
    defparam deldn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam deldn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO deldn_ibuf_preio (
            .PADOEN(N__6420),
            .PADOUT(N__6419),
            .PADIN(N__6418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(deldn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led2_obuf_iopad (
            .OE(N__6411),
            .DIN(N__6410),
            .DOUT(N__6409),
            .PACKAGEPIN(led2));
    defparam led2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led2_obuf_preio (
            .PADOEN(N__6411),
            .PADOUT(N__6410),
            .PADIN(N__6409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4811),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delup_ibuf_iopad (
            .OE(N__6402),
            .DIN(N__6401),
            .DOUT(N__6400),
            .PACKAGEPIN(delup));
    defparam delup_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delup_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delup_ibuf_preio (
            .PADOEN(N__6402),
            .PADOUT(N__6401),
            .PADIN(N__6400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delup_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led6_obuf_iopad (
            .OE(N__6393),
            .DIN(N__6392),
            .DOUT(N__6391),
            .PACKAGEPIN(led6));
    defparam led6_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led6_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led6_obuf_preio (
            .PADOEN(N__6393),
            .PADOUT(N__6392),
            .PADIN(N__6391),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3668),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led8_obuf_iopad (
            .OE(N__6384),
            .DIN(N__6383),
            .DOUT(N__6382),
            .PACKAGEPIN(led8));
    defparam led8_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led8_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led8_obuf_preio (
            .PADOEN(N__6384),
            .PADOUT(N__6383),
            .PADIN(N__6382),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3626),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led4_obuf_iopad (
            .OE(N__6375),
            .DIN(N__6374),
            .DOUT(N__6373),
            .PACKAGEPIN(led4));
    defparam led4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led4_obuf_preio (
            .PADOEN(N__6375),
            .PADOUT(N__6374),
            .PADIN(N__6373),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.io_0_iopad  (
            .OE(N__6366),
            .DIN(N__6365),
            .DOUT(N__6364),
            .PACKAGEPIN(apureset));
    defparam \arse.io_0_preio .PIN_TYPE=6'b010101;
    PRE_IO \arse.io_0_preio  (
            .PADOEN(N__6366),
            .PADOUT(N__6365),
            .PADIN(N__6364),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6080),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5914));
    IO_PAD lcol4_obuf_iopad (
            .OE(N__6357),
            .DIN(N__6356),
            .DOUT(N__6355),
            .PACKAGEPIN(lcol4));
    defparam lcol4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol4_obuf_preio (
            .PADOEN(N__6357),
            .PADOUT(N__6356),
            .PADIN(N__6355),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2540),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.diveight.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.diveight.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.diveight.io_0_iopad  (
            .OE(N__6348),
            .DIN(N__6347),
            .DOUT(N__6346),
            .PACKAGEPIN(cpuclk));
    defparam \arse.diveight.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.diveight.io_0_preio  (
            .PADOEN(N__6348),
            .PADOUT(N__6347),
            .PADIN(N__6346),
            .CLOCKENABLE(),
            .DOUT1(N__5975),
            .OUTPUTENABLE(N__4972),
            .DIN0(),
            .DOUT0(N__5804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5914));
    IO_PAD led5_obuf_iopad (
            .OE(N__6339),
            .DIN(N__6338),
            .DOUT(N__6337),
            .PACKAGEPIN(led5));
    defparam led5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led5_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led5_obuf_preio (
            .PADOEN(N__6339),
            .PADOUT(N__6338),
            .PADIN(N__6337),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4968),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD consolereset_ibuf_iopad (
            .OE(N__6330),
            .DIN(N__6329),
            .DOUT(N__6328),
            .PACKAGEPIN(consolereset));
    defparam consolereset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam consolereset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO consolereset_ibuf_preio (
            .PADOEN(N__6330),
            .PADOUT(N__6329),
            .PADIN(N__6328),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(consolereset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol2_obuf_iopad (
            .OE(N__6321),
            .DIN(N__6320),
            .DOUT(N__6319),
            .PACKAGEPIN(lcol2));
    defparam lcol2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol2_obuf_preio (
            .PADOEN(N__6321),
            .PADOUT(N__6320),
            .PADIN(N__6319),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3341),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led1_obuf_iopad (
            .OE(N__6312),
            .DIN(N__6311),
            .DOUT(N__6310),
            .PACKAGEPIN(led1));
    defparam led1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led1_obuf_preio (
            .PADOEN(N__6312),
            .PADOUT(N__6311),
            .PADIN(N__6310),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4949),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD apusync_ibuf_iopad (
            .OE(N__6303),
            .DIN(N__6302),
            .DOUT(N__6301),
            .PACKAGEPIN(apusync));
    defparam apusync_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam apusync_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO apusync_ibuf_preio (
            .PADOEN(N__6303),
            .PADOUT(N__6302),
            .PADIN(N__6301),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(apusync_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led7_obuf_iopad (
            .OE(N__6294),
            .DIN(N__6293),
            .DOUT(N__6292),
            .PACKAGEPIN(led7));
    defparam led7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led7_obuf_preio (
            .PADOEN(N__6294),
            .PADOUT(N__6293),
            .PADIN(N__6292),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3758),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol1_obuf_iopad (
            .OE(N__6285),
            .DIN(N__6284),
            .DOUT(N__6283),
            .PACKAGEPIN(lcol1));
    defparam lcol1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol1_obuf_preio (
            .PADOEN(N__6285),
            .PADOUT(N__6284),
            .PADIN(N__6283),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1505 (
            .O(N__6266),
            .I(N__6261));
    CascadeMux I__1504 (
            .O(N__6265),
            .I(N__6258));
    InMux I__1503 (
            .O(N__6264),
            .I(N__6252));
    InMux I__1502 (
            .O(N__6261),
            .I(N__6245));
    InMux I__1501 (
            .O(N__6258),
            .I(N__6245));
    InMux I__1500 (
            .O(N__6257),
            .I(N__6245));
    InMux I__1499 (
            .O(N__6256),
            .I(N__6240));
    InMux I__1498 (
            .O(N__6255),
            .I(N__6240));
    LocalMux I__1497 (
            .O(N__6252),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__1496 (
            .O(N__6245),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__1495 (
            .O(N__6240),
            .I(\arse.divseven.counterZ0Z_0 ));
    CascadeMux I__1494 (
            .O(N__6233),
            .I(N__6226));
    InMux I__1493 (
            .O(N__6232),
            .I(N__6222));
    InMux I__1492 (
            .O(N__6231),
            .I(N__6211));
    InMux I__1491 (
            .O(N__6230),
            .I(N__6211));
    InMux I__1490 (
            .O(N__6229),
            .I(N__6211));
    InMux I__1489 (
            .O(N__6226),
            .I(N__6211));
    InMux I__1488 (
            .O(N__6225),
            .I(N__6211));
    LocalMux I__1487 (
            .O(N__6222),
            .I(\arse.divseven.sevenZ0 ));
    LocalMux I__1486 (
            .O(N__6211),
            .I(\arse.divseven.sevenZ0 ));
    InMux I__1485 (
            .O(N__6206),
            .I(N__6203));
    LocalMux I__1484 (
            .O(N__6203),
            .I(N__6200));
    Span12Mux_v I__1483 (
            .O(N__6200),
            .I(N__6197));
    Odrv12 I__1482 (
            .O(N__6197),
            .I(apusync_c));
    CascadeMux I__1481 (
            .O(N__6194),
            .I(N__6191));
    InMux I__1480 (
            .O(N__6191),
            .I(N__6186));
    InMux I__1479 (
            .O(N__6190),
            .I(N__6183));
    InMux I__1478 (
            .O(N__6189),
            .I(N__6180));
    LocalMux I__1477 (
            .O(N__6186),
            .I(N__6175));
    LocalMux I__1476 (
            .O(N__6183),
            .I(N__6170));
    LocalMux I__1475 (
            .O(N__6180),
            .I(N__6170));
    InMux I__1474 (
            .O(N__6179),
            .I(N__6167));
    InMux I__1473 (
            .O(N__6178),
            .I(N__6164));
    Span4Mux_h I__1472 (
            .O(N__6175),
            .I(N__6157));
    Span4Mux_h I__1471 (
            .O(N__6170),
            .I(N__6157));
    LocalMux I__1470 (
            .O(N__6167),
            .I(N__6157));
    LocalMux I__1469 (
            .O(N__6164),
            .I(N__6154));
    Span4Mux_v I__1468 (
            .O(N__6157),
            .I(N__6148));
    Span4Mux_v I__1467 (
            .O(N__6154),
            .I(N__6148));
    InMux I__1466 (
            .O(N__6153),
            .I(N__6145));
    Odrv4 I__1465 (
            .O(N__6148),
            .I(\arse.apusynclatchedZ0 ));
    LocalMux I__1464 (
            .O(N__6145),
            .I(\arse.apusynclatchedZ0 ));
    InMux I__1463 (
            .O(N__6140),
            .I(N__6137));
    LocalMux I__1462 (
            .O(N__6137),
            .I(N__6134));
    Span4Mux_v I__1461 (
            .O(N__6134),
            .I(N__6129));
    InMux I__1460 (
            .O(N__6133),
            .I(N__6126));
    InMux I__1459 (
            .O(N__6132),
            .I(N__6123));
    Span4Mux_h I__1458 (
            .O(N__6129),
            .I(N__6120));
    LocalMux I__1457 (
            .O(N__6126),
            .I(N__6117));
    LocalMux I__1456 (
            .O(N__6123),
            .I(N__6114));
    Sp12to4 I__1455 (
            .O(N__6120),
            .I(N__6111));
    Span4Mux_v I__1454 (
            .O(N__6117),
            .I(N__6108));
    Span12Mux_s10_h I__1453 (
            .O(N__6114),
            .I(N__6104));
    Span12Mux_v I__1452 (
            .O(N__6111),
            .I(N__6099));
    Sp12to4 I__1451 (
            .O(N__6108),
            .I(N__6099));
    CascadeMux I__1450 (
            .O(N__6107),
            .I(N__6096));
    Span12Mux_v I__1449 (
            .O(N__6104),
            .I(N__6093));
    Span12Mux_h I__1448 (
            .O(N__6099),
            .I(N__6090));
    InMux I__1447 (
            .O(N__6096),
            .I(N__6087));
    Odrv12 I__1446 (
            .O(N__6093),
            .I(debouncedconsolereset));
    Odrv12 I__1445 (
            .O(N__6090),
            .I(debouncedconsolereset));
    LocalMux I__1444 (
            .O(N__6087),
            .I(debouncedconsolereset));
    IoInMux I__1443 (
            .O(N__6080),
            .I(N__6077));
    LocalMux I__1442 (
            .O(N__6077),
            .I(\arse.apuresetoutregZ0 ));
    InMux I__1441 (
            .O(N__6074),
            .I(N__6070));
    CascadeMux I__1440 (
            .O(N__6073),
            .I(N__6067));
    LocalMux I__1439 (
            .O(N__6070),
            .I(N__6062));
    InMux I__1438 (
            .O(N__6067),
            .I(N__6055));
    InMux I__1437 (
            .O(N__6066),
            .I(N__6055));
    InMux I__1436 (
            .O(N__6065),
            .I(N__6055));
    Odrv4 I__1435 (
            .O(N__6062),
            .I(\arse.diveight.counterZ0Z_0 ));
    LocalMux I__1434 (
            .O(N__6055),
            .I(\arse.diveight.counterZ0Z_0 ));
    InMux I__1433 (
            .O(N__6050),
            .I(N__6045));
    InMux I__1432 (
            .O(N__6049),
            .I(N__6042));
    InMux I__1431 (
            .O(N__6048),
            .I(N__6036));
    LocalMux I__1430 (
            .O(N__6045),
            .I(N__6031));
    LocalMux I__1429 (
            .O(N__6042),
            .I(N__6031));
    InMux I__1428 (
            .O(N__6041),
            .I(N__6024));
    InMux I__1427 (
            .O(N__6040),
            .I(N__6024));
    InMux I__1426 (
            .O(N__6039),
            .I(N__6024));
    LocalMux I__1425 (
            .O(N__6036),
            .I(\arse.cpuclkresetZ0 ));
    Odrv12 I__1424 (
            .O(N__6031),
            .I(\arse.cpuclkresetZ0 ));
    LocalMux I__1423 (
            .O(N__6024),
            .I(\arse.cpuclkresetZ0 ));
    CascadeMux I__1422 (
            .O(N__6017),
            .I(N__6014));
    InMux I__1421 (
            .O(N__6014),
            .I(N__6011));
    LocalMux I__1420 (
            .O(N__6011),
            .I(N__6006));
    InMux I__1419 (
            .O(N__6010),
            .I(N__6001));
    InMux I__1418 (
            .O(N__6009),
            .I(N__6001));
    Odrv4 I__1417 (
            .O(N__6006),
            .I(\arse.diveight.counterZ0Z_1 ));
    LocalMux I__1416 (
            .O(N__6001),
            .I(\arse.diveight.counterZ0Z_1 ));
    InMux I__1415 (
            .O(N__5996),
            .I(N__5993));
    LocalMux I__1414 (
            .O(N__5993),
            .I(N__5988));
    InMux I__1413 (
            .O(N__5992),
            .I(N__5985));
    InMux I__1412 (
            .O(N__5991),
            .I(N__5982));
    Odrv4 I__1411 (
            .O(N__5988),
            .I(\arse.diveight.counterZ0Z_2 ));
    LocalMux I__1410 (
            .O(N__5985),
            .I(\arse.diveight.counterZ0Z_2 ));
    LocalMux I__1409 (
            .O(N__5982),
            .I(\arse.diveight.counterZ0Z_2 ));
    IoInMux I__1408 (
            .O(N__5975),
            .I(N__5972));
    LocalMux I__1407 (
            .O(N__5972),
            .I(\arse.diveight.doutZ0Z_1 ));
    CascadeMux I__1406 (
            .O(N__5969),
            .I(N__5966));
    InMux I__1405 (
            .O(N__5966),
            .I(N__5963));
    LocalMux I__1404 (
            .O(N__5963),
            .I(\arse.divseven.N_46_0 ));
    CascadeMux I__1403 (
            .O(N__5960),
            .I(N__5955));
    CascadeMux I__1402 (
            .O(N__5959),
            .I(N__5949));
    InMux I__1401 (
            .O(N__5958),
            .I(N__5946));
    InMux I__1400 (
            .O(N__5955),
            .I(N__5939));
    InMux I__1399 (
            .O(N__5954),
            .I(N__5939));
    InMux I__1398 (
            .O(N__5953),
            .I(N__5939));
    InMux I__1397 (
            .O(N__5952),
            .I(N__5934));
    InMux I__1396 (
            .O(N__5949),
            .I(N__5934));
    LocalMux I__1395 (
            .O(N__5946),
            .I(\arse.divseven.counterZ0Z_1 ));
    LocalMux I__1394 (
            .O(N__5939),
            .I(\arse.divseven.counterZ0Z_1 ));
    LocalMux I__1393 (
            .O(N__5934),
            .I(\arse.divseven.counterZ0Z_1 ));
    InMux I__1392 (
            .O(N__5927),
            .I(N__5923));
    IoInMux I__1391 (
            .O(N__5926),
            .I(N__5920));
    LocalMux I__1390 (
            .O(N__5923),
            .I(\arse.divseven.doutZ0Z_1 ));
    LocalMux I__1389 (
            .O(N__5920),
            .I(\arse.divseven.doutZ0Z_1 ));
    ClkMux I__1388 (
            .O(N__5915),
            .I(N__5870));
    ClkMux I__1387 (
            .O(N__5914),
            .I(N__5870));
    ClkMux I__1386 (
            .O(N__5913),
            .I(N__5870));
    ClkMux I__1385 (
            .O(N__5912),
            .I(N__5870));
    ClkMux I__1384 (
            .O(N__5911),
            .I(N__5870));
    ClkMux I__1383 (
            .O(N__5910),
            .I(N__5870));
    ClkMux I__1382 (
            .O(N__5909),
            .I(N__5870));
    ClkMux I__1381 (
            .O(N__5908),
            .I(N__5870));
    ClkMux I__1380 (
            .O(N__5907),
            .I(N__5870));
    ClkMux I__1379 (
            .O(N__5906),
            .I(N__5870));
    ClkMux I__1378 (
            .O(N__5905),
            .I(N__5870));
    ClkMux I__1377 (
            .O(N__5904),
            .I(N__5870));
    ClkMux I__1376 (
            .O(N__5903),
            .I(N__5870));
    ClkMux I__1375 (
            .O(N__5902),
            .I(N__5870));
    ClkMux I__1374 (
            .O(N__5901),
            .I(N__5870));
    GlobalMux I__1373 (
            .O(N__5870),
            .I(N__5867));
    gio2CtrlBuf I__1372 (
            .O(N__5867),
            .I(PLLOUTCORE_g));
    InMux I__1371 (
            .O(N__5864),
            .I(N__5855));
    InMux I__1370 (
            .O(N__5863),
            .I(N__5852));
    InMux I__1369 (
            .O(N__5862),
            .I(N__5841));
    InMux I__1368 (
            .O(N__5861),
            .I(N__5841));
    InMux I__1367 (
            .O(N__5860),
            .I(N__5841));
    InMux I__1366 (
            .O(N__5859),
            .I(N__5841));
    InMux I__1365 (
            .O(N__5858),
            .I(N__5841));
    LocalMux I__1364 (
            .O(N__5855),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__1363 (
            .O(N__5852),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__1362 (
            .O(N__5841),
            .I(\arse.divseven.counterZ0Z_2 ));
    IoInMux I__1361 (
            .O(N__5834),
            .I(N__5831));
    LocalMux I__1360 (
            .O(N__5831),
            .I(\arse.divseven.doutZ0Z_0 ));
    CEMux I__1359 (
            .O(N__5828),
            .I(N__5825));
    LocalMux I__1358 (
            .O(N__5825),
            .I(N__5822));
    Odrv4 I__1357 (
            .O(N__5822),
            .I(\arse.divseven.un1_dout_2_sqmuxa_0_i ));
    CascadeMux I__1356 (
            .O(N__5819),
            .I(N__5815));
    InMux I__1355 (
            .O(N__5818),
            .I(N__5812));
    InMux I__1354 (
            .O(N__5815),
            .I(N__5809));
    LocalMux I__1353 (
            .O(N__5812),
            .I(\arse.doingsevenZ0 ));
    LocalMux I__1352 (
            .O(N__5809),
            .I(\arse.doingsevenZ0 ));
    IoInMux I__1351 (
            .O(N__5804),
            .I(N__5801));
    LocalMux I__1350 (
            .O(N__5801),
            .I(N__5798));
    Span4Mux_s0_h I__1349 (
            .O(N__5798),
            .I(N__5795));
    Odrv4 I__1348 (
            .O(N__5795),
            .I(\arse.diveight.doutZ1Z_0 ));
    InMux I__1347 (
            .O(N__5792),
            .I(N__5789));
    LocalMux I__1346 (
            .O(N__5789),
            .I(\arse.divseven.un1_counter_i_0_0 ));
    InMux I__1345 (
            .O(N__5786),
            .I(N__5781));
    InMux I__1344 (
            .O(N__5785),
            .I(N__5776));
    InMux I__1343 (
            .O(N__5784),
            .I(N__5773));
    LocalMux I__1342 (
            .O(N__5781),
            .I(N__5770));
    InMux I__1341 (
            .O(N__5780),
            .I(N__5765));
    InMux I__1340 (
            .O(N__5779),
            .I(N__5765));
    LocalMux I__1339 (
            .O(N__5776),
            .I(N__5760));
    LocalMux I__1338 (
            .O(N__5773),
            .I(N__5760));
    Span4Mux_h I__1337 (
            .O(N__5770),
            .I(N__5756));
    LocalMux I__1336 (
            .O(N__5765),
            .I(N__5751));
    Span4Mux_v I__1335 (
            .O(N__5760),
            .I(N__5751));
    InMux I__1334 (
            .O(N__5759),
            .I(N__5748));
    Span4Mux_h I__1333 (
            .O(N__5756),
            .I(N__5745));
    Odrv4 I__1332 (
            .O(N__5751),
            .I(delayConstantZ0Z_4));
    LocalMux I__1331 (
            .O(N__5748),
            .I(delayConstantZ0Z_4));
    Odrv4 I__1330 (
            .O(N__5745),
            .I(delayConstantZ0Z_4));
    InMux I__1329 (
            .O(N__5738),
            .I(N__5734));
    CascadeMux I__1328 (
            .O(N__5737),
            .I(N__5730));
    LocalMux I__1327 (
            .O(N__5734),
            .I(N__5725));
    InMux I__1326 (
            .O(N__5733),
            .I(N__5722));
    InMux I__1325 (
            .O(N__5730),
            .I(N__5719));
    InMux I__1324 (
            .O(N__5729),
            .I(N__5716));
    InMux I__1323 (
            .O(N__5728),
            .I(N__5713));
    Span4Mux_v I__1322 (
            .O(N__5725),
            .I(N__5709));
    LocalMux I__1321 (
            .O(N__5722),
            .I(N__5705));
    LocalMux I__1320 (
            .O(N__5719),
            .I(N__5698));
    LocalMux I__1319 (
            .O(N__5716),
            .I(N__5698));
    LocalMux I__1318 (
            .O(N__5713),
            .I(N__5698));
    InMux I__1317 (
            .O(N__5712),
            .I(N__5694));
    Sp12to4 I__1316 (
            .O(N__5709),
            .I(N__5691));
    InMux I__1315 (
            .O(N__5708),
            .I(N__5688));
    Span4Mux_v I__1314 (
            .O(N__5705),
            .I(N__5683));
    Span4Mux_v I__1313 (
            .O(N__5698),
            .I(N__5683));
    InMux I__1312 (
            .O(N__5697),
            .I(N__5680));
    LocalMux I__1311 (
            .O(N__5694),
            .I(delayConstantZ0Z_0));
    Odrv12 I__1310 (
            .O(N__5691),
            .I(delayConstantZ0Z_0));
    LocalMux I__1309 (
            .O(N__5688),
            .I(delayConstantZ0Z_0));
    Odrv4 I__1308 (
            .O(N__5683),
            .I(delayConstantZ0Z_0));
    LocalMux I__1307 (
            .O(N__5680),
            .I(delayConstantZ0Z_0));
    CascadeMux I__1306 (
            .O(N__5669),
            .I(N__5666));
    InMux I__1305 (
            .O(N__5666),
            .I(N__5663));
    LocalMux I__1304 (
            .O(N__5663),
            .I(N__5657));
    InMux I__1303 (
            .O(N__5662),
            .I(N__5654));
    InMux I__1302 (
            .O(N__5661),
            .I(N__5651));
    InMux I__1301 (
            .O(N__5660),
            .I(N__5648));
    Odrv4 I__1300 (
            .O(N__5657),
            .I(\arse.cpuresetcountZ0Z_0 ));
    LocalMux I__1299 (
            .O(N__5654),
            .I(\arse.cpuresetcountZ0Z_0 ));
    LocalMux I__1298 (
            .O(N__5651),
            .I(\arse.cpuresetcountZ0Z_0 ));
    LocalMux I__1297 (
            .O(N__5648),
            .I(\arse.cpuresetcountZ0Z_0 ));
    CascadeMux I__1296 (
            .O(N__5639),
            .I(N__5633));
    InMux I__1295 (
            .O(N__5638),
            .I(N__5630));
    InMux I__1294 (
            .O(N__5637),
            .I(N__5627));
    InMux I__1293 (
            .O(N__5636),
            .I(N__5624));
    InMux I__1292 (
            .O(N__5633),
            .I(N__5621));
    LocalMux I__1291 (
            .O(N__5630),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1290 (
            .O(N__5627),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1289 (
            .O(N__5624),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1288 (
            .O(N__5621),
            .I(\arse.cpuresetcountZ0Z_4 ));
    InMux I__1287 (
            .O(N__5612),
            .I(N__5609));
    LocalMux I__1286 (
            .O(N__5609),
            .I(\arse.g0_3 ));
    CascadeMux I__1285 (
            .O(N__5606),
            .I(\arse.g0_2_cascade_ ));
    InMux I__1284 (
            .O(N__5603),
            .I(N__5600));
    LocalMux I__1283 (
            .O(N__5600),
            .I(\arse.g0_4 ));
    InMux I__1282 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__1281 (
            .O(N__5594),
            .I(\arse.N_6 ));
    InMux I__1280 (
            .O(N__5591),
            .I(N__5588));
    LocalMux I__1279 (
            .O(N__5588),
            .I(\arse.g0_1 ));
    CascadeMux I__1278 (
            .O(N__5585),
            .I(\arse.g0_7_cascade_ ));
    CascadeMux I__1277 (
            .O(N__5582),
            .I(\arse.cpuresetoutreg_1_sqmuxa_cascade_ ));
    IoInMux I__1276 (
            .O(N__5579),
            .I(N__5576));
    LocalMux I__1275 (
            .O(N__5576),
            .I(N__5572));
    InMux I__1274 (
            .O(N__5575),
            .I(N__5569));
    Span4Mux_s3_h I__1273 (
            .O(N__5572),
            .I(N__5566));
    LocalMux I__1272 (
            .O(N__5569),
            .I(\arse.cpuresetoutregZ0 ));
    Odrv4 I__1271 (
            .O(N__5566),
            .I(\arse.cpuresetoutregZ0 ));
    InMux I__1270 (
            .O(N__5561),
            .I(N__5558));
    LocalMux I__1269 (
            .O(N__5558),
            .I(\arse.doingseven4 ));
    InMux I__1268 (
            .O(N__5555),
            .I(N__5552));
    LocalMux I__1267 (
            .O(N__5552),
            .I(\arse.doingseven3 ));
    SRMux I__1266 (
            .O(N__5549),
            .I(N__5544));
    SRMux I__1265 (
            .O(N__5548),
            .I(N__5541));
    SRMux I__1264 (
            .O(N__5547),
            .I(N__5537));
    LocalMux I__1263 (
            .O(N__5544),
            .I(N__5534));
    LocalMux I__1262 (
            .O(N__5541),
            .I(N__5531));
    SRMux I__1261 (
            .O(N__5540),
            .I(N__5528));
    LocalMux I__1260 (
            .O(N__5537),
            .I(N__5525));
    Odrv12 I__1259 (
            .O(N__5534),
            .I(debouncedconsolereset_i));
    Odrv12 I__1258 (
            .O(N__5531),
            .I(debouncedconsolereset_i));
    LocalMux I__1257 (
            .O(N__5528),
            .I(debouncedconsolereset_i));
    Odrv4 I__1256 (
            .O(N__5525),
            .I(debouncedconsolereset_i));
    InMux I__1255 (
            .O(N__5516),
            .I(\arse.un1_cpuresetcount_1_cry_6 ));
    CascadeMux I__1254 (
            .O(N__5513),
            .I(N__5509));
    CascadeMux I__1253 (
            .O(N__5512),
            .I(N__5503));
    InMux I__1252 (
            .O(N__5509),
            .I(N__5497));
    InMux I__1251 (
            .O(N__5508),
            .I(N__5497));
    InMux I__1250 (
            .O(N__5507),
            .I(N__5490));
    InMux I__1249 (
            .O(N__5506),
            .I(N__5486));
    InMux I__1248 (
            .O(N__5503),
            .I(N__5481));
    InMux I__1247 (
            .O(N__5502),
            .I(N__5481));
    LocalMux I__1246 (
            .O(N__5497),
            .I(N__5478));
    InMux I__1245 (
            .O(N__5496),
            .I(N__5473));
    InMux I__1244 (
            .O(N__5495),
            .I(N__5473));
    CascadeMux I__1243 (
            .O(N__5494),
            .I(N__5470));
    CascadeMux I__1242 (
            .O(N__5493),
            .I(N__5467));
    LocalMux I__1241 (
            .O(N__5490),
            .I(N__5463));
    InMux I__1240 (
            .O(N__5489),
            .I(N__5460));
    LocalMux I__1239 (
            .O(N__5486),
            .I(N__5457));
    LocalMux I__1238 (
            .O(N__5481),
            .I(N__5450));
    Span4Mux_h I__1237 (
            .O(N__5478),
            .I(N__5450));
    LocalMux I__1236 (
            .O(N__5473),
            .I(N__5450));
    InMux I__1235 (
            .O(N__5470),
            .I(N__5447));
    InMux I__1234 (
            .O(N__5467),
            .I(N__5442));
    InMux I__1233 (
            .O(N__5466),
            .I(N__5442));
    Span12Mux_s11_h I__1232 (
            .O(N__5463),
            .I(N__5437));
    LocalMux I__1231 (
            .O(N__5460),
            .I(N__5437));
    Span4Mux_v I__1230 (
            .O(N__5457),
            .I(N__5432));
    Span4Mux_v I__1229 (
            .O(N__5450),
            .I(N__5432));
    LocalMux I__1228 (
            .O(N__5447),
            .I(delayConstantZ0Z_1));
    LocalMux I__1227 (
            .O(N__5442),
            .I(delayConstantZ0Z_1));
    Odrv12 I__1226 (
            .O(N__5437),
            .I(delayConstantZ0Z_1));
    Odrv4 I__1225 (
            .O(N__5432),
            .I(delayConstantZ0Z_1));
    CascadeMux I__1224 (
            .O(N__5423),
            .I(N__5420));
    InMux I__1223 (
            .O(N__5420),
            .I(N__5411));
    CascadeMux I__1222 (
            .O(N__5419),
            .I(N__5408));
    CascadeMux I__1221 (
            .O(N__5418),
            .I(N__5402));
    CascadeMux I__1220 (
            .O(N__5417),
            .I(N__5399));
    CascadeMux I__1219 (
            .O(N__5416),
            .I(N__5396));
    CascadeMux I__1218 (
            .O(N__5415),
            .I(N__5393));
    CascadeMux I__1217 (
            .O(N__5414),
            .I(N__5390));
    LocalMux I__1216 (
            .O(N__5411),
            .I(N__5387));
    InMux I__1215 (
            .O(N__5408),
            .I(N__5382));
    CascadeMux I__1214 (
            .O(N__5407),
            .I(N__5379));
    CascadeMux I__1213 (
            .O(N__5406),
            .I(N__5376));
    InMux I__1212 (
            .O(N__5405),
            .I(N__5371));
    InMux I__1211 (
            .O(N__5402),
            .I(N__5371));
    InMux I__1210 (
            .O(N__5399),
            .I(N__5366));
    InMux I__1209 (
            .O(N__5396),
            .I(N__5366));
    InMux I__1208 (
            .O(N__5393),
            .I(N__5361));
    InMux I__1207 (
            .O(N__5390),
            .I(N__5361));
    Span4Mux_v I__1206 (
            .O(N__5387),
            .I(N__5358));
    CascadeMux I__1205 (
            .O(N__5386),
            .I(N__5355));
    InMux I__1204 (
            .O(N__5385),
            .I(N__5352));
    LocalMux I__1203 (
            .O(N__5382),
            .I(N__5349));
    InMux I__1202 (
            .O(N__5379),
            .I(N__5344));
    InMux I__1201 (
            .O(N__5376),
            .I(N__5344));
    LocalMux I__1200 (
            .O(N__5371),
            .I(N__5337));
    LocalMux I__1199 (
            .O(N__5366),
            .I(N__5337));
    LocalMux I__1198 (
            .O(N__5361),
            .I(N__5337));
    Sp12to4 I__1197 (
            .O(N__5358),
            .I(N__5334));
    InMux I__1196 (
            .O(N__5355),
            .I(N__5331));
    LocalMux I__1195 (
            .O(N__5352),
            .I(N__5322));
    Span4Mux_v I__1194 (
            .O(N__5349),
            .I(N__5322));
    LocalMux I__1193 (
            .O(N__5344),
            .I(N__5322));
    Span4Mux_v I__1192 (
            .O(N__5337),
            .I(N__5322));
    Odrv12 I__1191 (
            .O(N__5334),
            .I(delayConstantZ0Z_5));
    LocalMux I__1190 (
            .O(N__5331),
            .I(delayConstantZ0Z_5));
    Odrv4 I__1189 (
            .O(N__5322),
            .I(delayConstantZ0Z_5));
    InMux I__1188 (
            .O(N__5315),
            .I(N__5312));
    LocalMux I__1187 (
            .O(N__5312),
            .I(\arse.g0_i_a3_4 ));
    InMux I__1186 (
            .O(N__5309),
            .I(N__5303));
    InMux I__1185 (
            .O(N__5308),
            .I(N__5300));
    InMux I__1184 (
            .O(N__5307),
            .I(N__5297));
    InMux I__1183 (
            .O(N__5306),
            .I(N__5294));
    LocalMux I__1182 (
            .O(N__5303),
            .I(\arse.cpuresetcountZ0Z_5 ));
    LocalMux I__1181 (
            .O(N__5300),
            .I(\arse.cpuresetcountZ0Z_5 ));
    LocalMux I__1180 (
            .O(N__5297),
            .I(\arse.cpuresetcountZ0Z_5 ));
    LocalMux I__1179 (
            .O(N__5294),
            .I(\arse.cpuresetcountZ0Z_5 ));
    CascadeMux I__1178 (
            .O(N__5285),
            .I(\arse.doingseven3_6_cascade_ ));
    InMux I__1177 (
            .O(N__5282),
            .I(N__5276));
    InMux I__1176 (
            .O(N__5281),
            .I(N__5273));
    InMux I__1175 (
            .O(N__5280),
            .I(N__5270));
    InMux I__1174 (
            .O(N__5279),
            .I(N__5267));
    LocalMux I__1173 (
            .O(N__5276),
            .I(\arse.cpuresetcountZ0Z_1 ));
    LocalMux I__1172 (
            .O(N__5273),
            .I(\arse.cpuresetcountZ0Z_1 ));
    LocalMux I__1171 (
            .O(N__5270),
            .I(\arse.cpuresetcountZ0Z_1 ));
    LocalMux I__1170 (
            .O(N__5267),
            .I(\arse.cpuresetcountZ0Z_1 ));
    InMux I__1169 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__1168 (
            .O(N__5255),
            .I(\arse.doingseven3_1 ));
    InMux I__1167 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__1166 (
            .O(N__5249),
            .I(\arse.doingseven3_6 ));
    CascadeMux I__1165 (
            .O(N__5246),
            .I(\arse.doingseven3_1_cascade_ ));
    InMux I__1164 (
            .O(N__5243),
            .I(N__5240));
    LocalMux I__1163 (
            .O(N__5240),
            .I(N__5237));
    Span4Mux_v I__1162 (
            .O(N__5237),
            .I(N__5234));
    Span4Mux_h I__1161 (
            .O(N__5234),
            .I(N__5231));
    Odrv4 I__1160 (
            .O(N__5231),
            .I(delayConstant_fastZ0Z_6));
    InMux I__1159 (
            .O(N__5228),
            .I(N__5225));
    LocalMux I__1158 (
            .O(N__5225),
            .I(N__5222));
    Span4Mux_h I__1157 (
            .O(N__5222),
            .I(N__5219));
    Span4Mux_h I__1156 (
            .O(N__5219),
            .I(N__5216));
    Odrv4 I__1155 (
            .O(N__5216),
            .I(delayConstant_fastZ0Z_2));
    CascadeMux I__1154 (
            .O(N__5213),
            .I(N__5207));
    CascadeMux I__1153 (
            .O(N__5212),
            .I(N__5204));
    CascadeMux I__1152 (
            .O(N__5211),
            .I(N__5201));
    InMux I__1151 (
            .O(N__5210),
            .I(N__5198));
    InMux I__1150 (
            .O(N__5207),
            .I(N__5195));
    InMux I__1149 (
            .O(N__5204),
            .I(N__5190));
    InMux I__1148 (
            .O(N__5201),
            .I(N__5190));
    LocalMux I__1147 (
            .O(N__5198),
            .I(\arse.cpuresetcountZ0Z_6 ));
    LocalMux I__1146 (
            .O(N__5195),
            .I(\arse.cpuresetcountZ0Z_6 ));
    LocalMux I__1145 (
            .O(N__5190),
            .I(\arse.cpuresetcountZ0Z_6 ));
    InMux I__1144 (
            .O(N__5183),
            .I(N__5175));
    InMux I__1143 (
            .O(N__5182),
            .I(N__5175));
    InMux I__1142 (
            .O(N__5181),
            .I(N__5172));
    InMux I__1141 (
            .O(N__5180),
            .I(N__5169));
    LocalMux I__1140 (
            .O(N__5175),
            .I(\arse.cpuresetcountZ0Z_2 ));
    LocalMux I__1139 (
            .O(N__5172),
            .I(\arse.cpuresetcountZ0Z_2 ));
    LocalMux I__1138 (
            .O(N__5169),
            .I(\arse.cpuresetcountZ0Z_2 ));
    InMux I__1137 (
            .O(N__5162),
            .I(N__5159));
    LocalMux I__1136 (
            .O(N__5159),
            .I(N__5155));
    CascadeMux I__1135 (
            .O(N__5158),
            .I(N__5148));
    Span4Mux_h I__1134 (
            .O(N__5155),
            .I(N__5144));
    InMux I__1133 (
            .O(N__5154),
            .I(N__5141));
    CascadeMux I__1132 (
            .O(N__5153),
            .I(N__5138));
    InMux I__1131 (
            .O(N__5152),
            .I(N__5135));
    InMux I__1130 (
            .O(N__5151),
            .I(N__5132));
    InMux I__1129 (
            .O(N__5148),
            .I(N__5129));
    InMux I__1128 (
            .O(N__5147),
            .I(N__5126));
    Span4Mux_v I__1127 (
            .O(N__5144),
            .I(N__5123));
    LocalMux I__1126 (
            .O(N__5141),
            .I(N__5120));
    InMux I__1125 (
            .O(N__5138),
            .I(N__5117));
    LocalMux I__1124 (
            .O(N__5135),
            .I(N__5112));
    LocalMux I__1123 (
            .O(N__5132),
            .I(N__5112));
    LocalMux I__1122 (
            .O(N__5129),
            .I(N__5107));
    LocalMux I__1121 (
            .O(N__5126),
            .I(N__5107));
    Span4Mux_h I__1120 (
            .O(N__5123),
            .I(N__5102));
    Span4Mux_v I__1119 (
            .O(N__5120),
            .I(N__5102));
    LocalMux I__1118 (
            .O(N__5117),
            .I(delayConstantZ0Z_7));
    Odrv12 I__1117 (
            .O(N__5112),
            .I(delayConstantZ0Z_7));
    Odrv4 I__1116 (
            .O(N__5107),
            .I(delayConstantZ0Z_7));
    Odrv4 I__1115 (
            .O(N__5102),
            .I(delayConstantZ0Z_7));
    InMux I__1114 (
            .O(N__5093),
            .I(N__5089));
    CascadeMux I__1113 (
            .O(N__5092),
            .I(N__5084));
    LocalMux I__1112 (
            .O(N__5089),
            .I(N__5079));
    InMux I__1111 (
            .O(N__5088),
            .I(N__5076));
    InMux I__1110 (
            .O(N__5087),
            .I(N__5073));
    InMux I__1109 (
            .O(N__5084),
            .I(N__5070));
    InMux I__1108 (
            .O(N__5083),
            .I(N__5065));
    InMux I__1107 (
            .O(N__5082),
            .I(N__5065));
    Span4Mux_h I__1106 (
            .O(N__5079),
            .I(N__5062));
    LocalMux I__1105 (
            .O(N__5076),
            .I(N__5059));
    LocalMux I__1104 (
            .O(N__5073),
            .I(N__5055));
    LocalMux I__1103 (
            .O(N__5070),
            .I(N__5052));
    LocalMux I__1102 (
            .O(N__5065),
            .I(N__5049));
    Span4Mux_v I__1101 (
            .O(N__5062),
            .I(N__5046));
    Span4Mux_h I__1100 (
            .O(N__5059),
            .I(N__5043));
    InMux I__1099 (
            .O(N__5058),
            .I(N__5040));
    Span4Mux_h I__1098 (
            .O(N__5055),
            .I(N__5037));
    Span4Mux_v I__1097 (
            .O(N__5052),
            .I(N__5032));
    Span4Mux_v I__1096 (
            .O(N__5049),
            .I(N__5032));
    Odrv4 I__1095 (
            .O(N__5046),
            .I(delayConstantZ0Z_3));
    Odrv4 I__1094 (
            .O(N__5043),
            .I(delayConstantZ0Z_3));
    LocalMux I__1093 (
            .O(N__5040),
            .I(delayConstantZ0Z_3));
    Odrv4 I__1092 (
            .O(N__5037),
            .I(delayConstantZ0Z_3));
    Odrv4 I__1091 (
            .O(N__5032),
            .I(delayConstantZ0Z_3));
    CascadeMux I__1090 (
            .O(N__5021),
            .I(N__5017));
    InMux I__1089 (
            .O(N__5020),
            .I(N__5012));
    InMux I__1088 (
            .O(N__5017),
            .I(N__5009));
    InMux I__1087 (
            .O(N__5016),
            .I(N__5004));
    InMux I__1086 (
            .O(N__5015),
            .I(N__5004));
    LocalMux I__1085 (
            .O(N__5012),
            .I(\arse.cpuresetcountZ0Z_7 ));
    LocalMux I__1084 (
            .O(N__5009),
            .I(\arse.cpuresetcountZ0Z_7 ));
    LocalMux I__1083 (
            .O(N__5004),
            .I(\arse.cpuresetcountZ0Z_7 ));
    InMux I__1082 (
            .O(N__4997),
            .I(N__4990));
    InMux I__1081 (
            .O(N__4996),
            .I(N__4983));
    InMux I__1080 (
            .O(N__4995),
            .I(N__4983));
    InMux I__1079 (
            .O(N__4994),
            .I(N__4983));
    InMux I__1078 (
            .O(N__4993),
            .I(N__4980));
    LocalMux I__1077 (
            .O(N__4990),
            .I(\arse.cpuresetcountZ0Z_3 ));
    LocalMux I__1076 (
            .O(N__4983),
            .I(\arse.cpuresetcountZ0Z_3 ));
    LocalMux I__1075 (
            .O(N__4980),
            .I(\arse.cpuresetcountZ0Z_3 ));
    IoInMux I__1074 (
            .O(N__4973),
            .I(N__4969));
    IoInMux I__1073 (
            .O(N__4972),
            .I(N__4965));
    LocalMux I__1072 (
            .O(N__4969),
            .I(N__4962));
    IoInMux I__1071 (
            .O(N__4968),
            .I(N__4959));
    LocalMux I__1070 (
            .O(N__4965),
            .I(N__4956));
    Span4Mux_s3_h I__1069 (
            .O(N__4962),
            .I(N__4953));
    LocalMux I__1068 (
            .O(N__4959),
            .I(N__4950));
    IoSpan4Mux I__1067 (
            .O(N__4956),
            .I(N__4946));
    Span4Mux_v I__1066 (
            .O(N__4953),
            .I(N__4943));
    IoSpan4Mux I__1065 (
            .O(N__4950),
            .I(N__4940));
    IoInMux I__1064 (
            .O(N__4949),
            .I(N__4937));
    Sp12to4 I__1063 (
            .O(N__4946),
            .I(N__4934));
    Sp12to4 I__1062 (
            .O(N__4943),
            .I(N__4931));
    IoSpan4Mux I__1061 (
            .O(N__4940),
            .I(N__4928));
    LocalMux I__1060 (
            .O(N__4937),
            .I(N__4925));
    Span12Mux_s9_h I__1059 (
            .O(N__4934),
            .I(N__4922));
    Span12Mux_s9_h I__1058 (
            .O(N__4931),
            .I(N__4919));
    Span4Mux_s1_v I__1057 (
            .O(N__4928),
            .I(N__4914));
    Span4Mux_s1_v I__1056 (
            .O(N__4925),
            .I(N__4914));
    Span12Mux_v I__1055 (
            .O(N__4922),
            .I(N__4911));
    Span12Mux_v I__1054 (
            .O(N__4919),
            .I(N__4908));
    Span4Mux_v I__1053 (
            .O(N__4914),
            .I(N__4905));
    Odrv12 I__1052 (
            .O(N__4911),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1051 (
            .O(N__4908),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1050 (
            .O(N__4905),
            .I(CONSTANT_ONE_NET));
    InMux I__1049 (
            .O(N__4898),
            .I(\arse.un1_cpuresetcount_1_cry_0 ));
    InMux I__1048 (
            .O(N__4895),
            .I(\arse.un1_cpuresetcount_1_cry_1 ));
    InMux I__1047 (
            .O(N__4892),
            .I(\arse.un1_cpuresetcount_1_cry_2 ));
    InMux I__1046 (
            .O(N__4889),
            .I(\arse.un1_cpuresetcount_1_cry_3 ));
    InMux I__1045 (
            .O(N__4886),
            .I(\arse.un1_cpuresetcount_1_cry_4 ));
    InMux I__1044 (
            .O(N__4883),
            .I(\arse.un1_cpuresetcount_1_cry_5 ));
    InMux I__1043 (
            .O(N__4880),
            .I(N__4877));
    LocalMux I__1042 (
            .O(N__4877),
            .I(\dig1.N_25 ));
    CascadeMux I__1041 (
            .O(N__4874),
            .I(\dig1.N_22_cascade_ ));
    InMux I__1040 (
            .O(N__4871),
            .I(N__4868));
    LocalMux I__1039 (
            .O(N__4868),
            .I(\dig1.leds_17_i_0_ns_1_2 ));
    InMux I__1038 (
            .O(N__4865),
            .I(N__4861));
    InMux I__1037 (
            .O(N__4864),
            .I(N__4858));
    LocalMux I__1036 (
            .O(N__4861),
            .I(un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2));
    LocalMux I__1035 (
            .O(N__4858),
            .I(un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2));
    InMux I__1034 (
            .O(N__4853),
            .I(N__4849));
    InMux I__1033 (
            .O(N__4852),
            .I(N__4846));
    LocalMux I__1032 (
            .O(N__4849),
            .I(un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92));
    LocalMux I__1031 (
            .O(N__4846),
            .I(un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92));
    SRMux I__1030 (
            .O(N__4841),
            .I(N__4817));
    SRMux I__1029 (
            .O(N__4840),
            .I(N__4817));
    SRMux I__1028 (
            .O(N__4839),
            .I(N__4817));
    SRMux I__1027 (
            .O(N__4838),
            .I(N__4817));
    SRMux I__1026 (
            .O(N__4837),
            .I(N__4817));
    SRMux I__1025 (
            .O(N__4836),
            .I(N__4817));
    SRMux I__1024 (
            .O(N__4835),
            .I(N__4817));
    SRMux I__1023 (
            .O(N__4834),
            .I(N__4817));
    GlobalMux I__1022 (
            .O(N__4817),
            .I(N__4814));
    gio2CtrlBuf I__1021 (
            .O(N__4814),
            .I(masterreset_c_i_g));
    IoInMux I__1020 (
            .O(N__4811),
            .I(N__4808));
    LocalMux I__1019 (
            .O(N__4808),
            .I(N__4805));
    IoSpan4Mux I__1018 (
            .O(N__4805),
            .I(N__4802));
    Span4Mux_s3_v I__1017 (
            .O(N__4802),
            .I(N__4799));
    Sp12to4 I__1016 (
            .O(N__4799),
            .I(N__4796));
    Span12Mux_s11_v I__1015 (
            .O(N__4796),
            .I(N__4793));
    Odrv12 I__1014 (
            .O(N__4793),
            .I(leds_1_i_0_1));
    InMux I__1013 (
            .O(N__4790),
            .I(N__4787));
    LocalMux I__1012 (
            .O(N__4787),
            .I(N__4757));
    ClkMux I__1011 (
            .O(N__4786),
            .I(N__4700));
    ClkMux I__1010 (
            .O(N__4785),
            .I(N__4700));
    ClkMux I__1009 (
            .O(N__4784),
            .I(N__4700));
    ClkMux I__1008 (
            .O(N__4783),
            .I(N__4700));
    ClkMux I__1007 (
            .O(N__4782),
            .I(N__4700));
    ClkMux I__1006 (
            .O(N__4781),
            .I(N__4700));
    ClkMux I__1005 (
            .O(N__4780),
            .I(N__4700));
    ClkMux I__1004 (
            .O(N__4779),
            .I(N__4700));
    ClkMux I__1003 (
            .O(N__4778),
            .I(N__4700));
    ClkMux I__1002 (
            .O(N__4777),
            .I(N__4700));
    ClkMux I__1001 (
            .O(N__4776),
            .I(N__4700));
    ClkMux I__1000 (
            .O(N__4775),
            .I(N__4700));
    ClkMux I__999 (
            .O(N__4774),
            .I(N__4700));
    ClkMux I__998 (
            .O(N__4773),
            .I(N__4700));
    ClkMux I__997 (
            .O(N__4772),
            .I(N__4700));
    ClkMux I__996 (
            .O(N__4771),
            .I(N__4700));
    ClkMux I__995 (
            .O(N__4770),
            .I(N__4700));
    ClkMux I__994 (
            .O(N__4769),
            .I(N__4700));
    ClkMux I__993 (
            .O(N__4768),
            .I(N__4700));
    ClkMux I__992 (
            .O(N__4767),
            .I(N__4700));
    ClkMux I__991 (
            .O(N__4766),
            .I(N__4700));
    ClkMux I__990 (
            .O(N__4765),
            .I(N__4700));
    ClkMux I__989 (
            .O(N__4764),
            .I(N__4700));
    ClkMux I__988 (
            .O(N__4763),
            .I(N__4700));
    ClkMux I__987 (
            .O(N__4762),
            .I(N__4700));
    ClkMux I__986 (
            .O(N__4761),
            .I(N__4700));
    ClkMux I__985 (
            .O(N__4760),
            .I(N__4700));
    Glb2LocalMux I__984 (
            .O(N__4757),
            .I(N__4700));
    GlobalMux I__983 (
            .O(N__4700),
            .I(N__4697));
    gio2CtrlBuf I__982 (
            .O(N__4697),
            .I(PACKAGEPIN_0_c_g));
    CEMux I__981 (
            .O(N__4694),
            .I(N__4691));
    LocalMux I__980 (
            .O(N__4691),
            .I(N__4686));
    CEMux I__979 (
            .O(N__4690),
            .I(N__4683));
    CEMux I__978 (
            .O(N__4689),
            .I(N__4675));
    Span4Mux_v I__977 (
            .O(N__4686),
            .I(N__4670));
    LocalMux I__976 (
            .O(N__4683),
            .I(N__4670));
    CEMux I__975 (
            .O(N__4682),
            .I(N__4667));
    CEMux I__974 (
            .O(N__4681),
            .I(N__4657));
    CEMux I__973 (
            .O(N__4680),
            .I(N__4654));
    InMux I__972 (
            .O(N__4679),
            .I(N__4651));
    InMux I__971 (
            .O(N__4678),
            .I(N__4648));
    LocalMux I__970 (
            .O(N__4675),
            .I(N__4645));
    Span4Mux_h I__969 (
            .O(N__4670),
            .I(N__4640));
    LocalMux I__968 (
            .O(N__4667),
            .I(N__4640));
    CascadeMux I__967 (
            .O(N__4666),
            .I(N__4634));
    CascadeMux I__966 (
            .O(N__4665),
            .I(N__4630));
    CascadeMux I__965 (
            .O(N__4664),
            .I(N__4626));
    CascadeMux I__964 (
            .O(N__4663),
            .I(N__4623));
    CascadeMux I__963 (
            .O(N__4662),
            .I(N__4620));
    CEMux I__962 (
            .O(N__4661),
            .I(N__4614));
    InMux I__961 (
            .O(N__4660),
            .I(N__4611));
    LocalMux I__960 (
            .O(N__4657),
            .I(N__4606));
    LocalMux I__959 (
            .O(N__4654),
            .I(N__4606));
    LocalMux I__958 (
            .O(N__4651),
            .I(N__4601));
    LocalMux I__957 (
            .O(N__4648),
            .I(N__4601));
    Span4Mux_v I__956 (
            .O(N__4645),
            .I(N__4596));
    Span4Mux_h I__955 (
            .O(N__4640),
            .I(N__4596));
    CascadeMux I__954 (
            .O(N__4639),
            .I(N__4592));
    CascadeMux I__953 (
            .O(N__4638),
            .I(N__4589));
    InMux I__952 (
            .O(N__4637),
            .I(N__4583));
    InMux I__951 (
            .O(N__4634),
            .I(N__4580));
    InMux I__950 (
            .O(N__4633),
            .I(N__4577));
    InMux I__949 (
            .O(N__4630),
            .I(N__4572));
    InMux I__948 (
            .O(N__4629),
            .I(N__4572));
    InMux I__947 (
            .O(N__4626),
            .I(N__4569));
    InMux I__946 (
            .O(N__4623),
            .I(N__4564));
    InMux I__945 (
            .O(N__4620),
            .I(N__4564));
    InMux I__944 (
            .O(N__4619),
            .I(N__4557));
    InMux I__943 (
            .O(N__4618),
            .I(N__4557));
    InMux I__942 (
            .O(N__4617),
            .I(N__4557));
    LocalMux I__941 (
            .O(N__4614),
            .I(N__4554));
    LocalMux I__940 (
            .O(N__4611),
            .I(N__4549));
    Span4Mux_v I__939 (
            .O(N__4606),
            .I(N__4549));
    Span4Mux_h I__938 (
            .O(N__4601),
            .I(N__4544));
    Span4Mux_h I__937 (
            .O(N__4596),
            .I(N__4544));
    InMux I__936 (
            .O(N__4595),
            .I(N__4539));
    InMux I__935 (
            .O(N__4592),
            .I(N__4539));
    InMux I__934 (
            .O(N__4589),
            .I(N__4530));
    InMux I__933 (
            .O(N__4588),
            .I(N__4530));
    InMux I__932 (
            .O(N__4587),
            .I(N__4530));
    InMux I__931 (
            .O(N__4586),
            .I(N__4530));
    LocalMux I__930 (
            .O(N__4583),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__929 (
            .O(N__4580),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__928 (
            .O(N__4577),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__927 (
            .O(N__4572),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__926 (
            .O(N__4569),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__925 (
            .O(N__4564),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__924 (
            .O(N__4557),
            .I(clock_out_RNIR6ER_0));
    Odrv12 I__923 (
            .O(N__4554),
            .I(clock_out_RNIR6ER_0));
    Odrv4 I__922 (
            .O(N__4549),
            .I(clock_out_RNIR6ER_0));
    Odrv4 I__921 (
            .O(N__4544),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__920 (
            .O(N__4539),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__919 (
            .O(N__4530),
            .I(clock_out_RNIR6ER_0));
    CascadeMux I__918 (
            .O(N__4505),
            .I(\dig1.N_52_cascade_ ));
    InMux I__917 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__916 (
            .O(N__4499),
            .I(\dig1.N_54 ));
    InMux I__915 (
            .O(N__4496),
            .I(N__4493));
    LocalMux I__914 (
            .O(N__4493),
            .I(\dig1.N_55 ));
    CascadeMux I__913 (
            .O(N__4490),
            .I(N__4485));
    InMux I__912 (
            .O(N__4489),
            .I(N__4480));
    InMux I__911 (
            .O(N__4488),
            .I(N__4480));
    InMux I__910 (
            .O(N__4485),
            .I(N__4477));
    LocalMux I__909 (
            .O(N__4480),
            .I(N__4467));
    LocalMux I__908 (
            .O(N__4477),
            .I(N__4460));
    InMux I__907 (
            .O(N__4476),
            .I(N__4455));
    InMux I__906 (
            .O(N__4475),
            .I(N__4455));
    InMux I__905 (
            .O(N__4474),
            .I(N__4440));
    InMux I__904 (
            .O(N__4473),
            .I(N__4435));
    InMux I__903 (
            .O(N__4472),
            .I(N__4435));
    InMux I__902 (
            .O(N__4471),
            .I(N__4432));
    InMux I__901 (
            .O(N__4470),
            .I(N__4429));
    Span4Mux_h I__900 (
            .O(N__4467),
            .I(N__4426));
    InMux I__899 (
            .O(N__4466),
            .I(N__4421));
    InMux I__898 (
            .O(N__4465),
            .I(N__4421));
    InMux I__897 (
            .O(N__4464),
            .I(N__4416));
    InMux I__896 (
            .O(N__4463),
            .I(N__4416));
    Span4Mux_v I__895 (
            .O(N__4460),
            .I(N__4411));
    LocalMux I__894 (
            .O(N__4455),
            .I(N__4411));
    InMux I__893 (
            .O(N__4454),
            .I(N__4406));
    InMux I__892 (
            .O(N__4453),
            .I(N__4406));
    InMux I__891 (
            .O(N__4452),
            .I(N__4401));
    InMux I__890 (
            .O(N__4451),
            .I(N__4401));
    InMux I__889 (
            .O(N__4450),
            .I(N__4394));
    InMux I__888 (
            .O(N__4449),
            .I(N__4394));
    InMux I__887 (
            .O(N__4448),
            .I(N__4394));
    InMux I__886 (
            .O(N__4447),
            .I(N__4389));
    InMux I__885 (
            .O(N__4446),
            .I(N__4389));
    InMux I__884 (
            .O(N__4445),
            .I(N__4382));
    InMux I__883 (
            .O(N__4444),
            .I(N__4382));
    InMux I__882 (
            .O(N__4443),
            .I(N__4382));
    LocalMux I__881 (
            .O(N__4440),
            .I(N__4377));
    LocalMux I__880 (
            .O(N__4435),
            .I(N__4377));
    LocalMux I__879 (
            .O(N__4432),
            .I(colZ0Z_0));
    LocalMux I__878 (
            .O(N__4429),
            .I(colZ0Z_0));
    Odrv4 I__877 (
            .O(N__4426),
            .I(colZ0Z_0));
    LocalMux I__876 (
            .O(N__4421),
            .I(colZ0Z_0));
    LocalMux I__875 (
            .O(N__4416),
            .I(colZ0Z_0));
    Odrv4 I__874 (
            .O(N__4411),
            .I(colZ0Z_0));
    LocalMux I__873 (
            .O(N__4406),
            .I(colZ0Z_0));
    LocalMux I__872 (
            .O(N__4401),
            .I(colZ0Z_0));
    LocalMux I__871 (
            .O(N__4394),
            .I(colZ0Z_0));
    LocalMux I__870 (
            .O(N__4389),
            .I(colZ0Z_0));
    LocalMux I__869 (
            .O(N__4382),
            .I(colZ0Z_0));
    Odrv12 I__868 (
            .O(N__4377),
            .I(colZ0Z_0));
    InMux I__867 (
            .O(N__4352),
            .I(N__4344));
    InMux I__866 (
            .O(N__4351),
            .I(N__4344));
    CascadeMux I__865 (
            .O(N__4350),
            .I(N__4341));
    InMux I__864 (
            .O(N__4349),
            .I(N__4338));
    LocalMux I__863 (
            .O(N__4344),
            .I(N__4326));
    InMux I__862 (
            .O(N__4341),
            .I(N__4323));
    LocalMux I__861 (
            .O(N__4338),
            .I(N__4319));
    InMux I__860 (
            .O(N__4337),
            .I(N__4314));
    InMux I__859 (
            .O(N__4336),
            .I(N__4314));
    InMux I__858 (
            .O(N__4335),
            .I(N__4301));
    InMux I__857 (
            .O(N__4334),
            .I(N__4296));
    InMux I__856 (
            .O(N__4333),
            .I(N__4296));
    InMux I__855 (
            .O(N__4332),
            .I(N__4291));
    InMux I__854 (
            .O(N__4331),
            .I(N__4291));
    InMux I__853 (
            .O(N__4330),
            .I(N__4288));
    InMux I__852 (
            .O(N__4329),
            .I(N__4285));
    Span4Mux_h I__851 (
            .O(N__4326),
            .I(N__4282));
    LocalMux I__850 (
            .O(N__4323),
            .I(N__4279));
    InMux I__849 (
            .O(N__4322),
            .I(N__4276));
    Span4Mux_v I__848 (
            .O(N__4319),
            .I(N__4271));
    LocalMux I__847 (
            .O(N__4314),
            .I(N__4271));
    InMux I__846 (
            .O(N__4313),
            .I(N__4266));
    InMux I__845 (
            .O(N__4312),
            .I(N__4266));
    InMux I__844 (
            .O(N__4311),
            .I(N__4259));
    InMux I__843 (
            .O(N__4310),
            .I(N__4259));
    InMux I__842 (
            .O(N__4309),
            .I(N__4259));
    InMux I__841 (
            .O(N__4308),
            .I(N__4254));
    InMux I__840 (
            .O(N__4307),
            .I(N__4254));
    InMux I__839 (
            .O(N__4306),
            .I(N__4247));
    InMux I__838 (
            .O(N__4305),
            .I(N__4247));
    InMux I__837 (
            .O(N__4304),
            .I(N__4247));
    LocalMux I__836 (
            .O(N__4301),
            .I(N__4240));
    LocalMux I__835 (
            .O(N__4296),
            .I(N__4240));
    LocalMux I__834 (
            .O(N__4291),
            .I(N__4240));
    LocalMux I__833 (
            .O(N__4288),
            .I(colZ0Z_1));
    LocalMux I__832 (
            .O(N__4285),
            .I(colZ0Z_1));
    Odrv4 I__831 (
            .O(N__4282),
            .I(colZ0Z_1));
    Odrv4 I__830 (
            .O(N__4279),
            .I(colZ0Z_1));
    LocalMux I__829 (
            .O(N__4276),
            .I(colZ0Z_1));
    Odrv4 I__828 (
            .O(N__4271),
            .I(colZ0Z_1));
    LocalMux I__827 (
            .O(N__4266),
            .I(colZ0Z_1));
    LocalMux I__826 (
            .O(N__4259),
            .I(colZ0Z_1));
    LocalMux I__825 (
            .O(N__4254),
            .I(colZ0Z_1));
    LocalMux I__824 (
            .O(N__4247),
            .I(colZ0Z_1));
    Odrv4 I__823 (
            .O(N__4240),
            .I(colZ0Z_1));
    CascadeMux I__822 (
            .O(N__4217),
            .I(N__4209));
    CascadeMux I__821 (
            .O(N__4216),
            .I(N__4205));
    CascadeMux I__820 (
            .O(N__4215),
            .I(N__4202));
    CascadeMux I__819 (
            .O(N__4214),
            .I(N__4198));
    CascadeMux I__818 (
            .O(N__4213),
            .I(N__4192));
    InMux I__817 (
            .O(N__4212),
            .I(N__4187));
    InMux I__816 (
            .O(N__4209),
            .I(N__4187));
    CascadeMux I__815 (
            .O(N__4208),
            .I(N__4184));
    InMux I__814 (
            .O(N__4205),
            .I(N__4179));
    InMux I__813 (
            .O(N__4202),
            .I(N__4179));
    InMux I__812 (
            .O(N__4201),
            .I(N__4176));
    InMux I__811 (
            .O(N__4198),
            .I(N__4173));
    CascadeMux I__810 (
            .O(N__4197),
            .I(N__4169));
    InMux I__809 (
            .O(N__4196),
            .I(N__4166));
    InMux I__808 (
            .O(N__4195),
            .I(N__4161));
    InMux I__807 (
            .O(N__4192),
            .I(N__4161));
    LocalMux I__806 (
            .O(N__4187),
            .I(N__4158));
    InMux I__805 (
            .O(N__4184),
            .I(N__4155));
    LocalMux I__804 (
            .O(N__4179),
            .I(N__4152));
    LocalMux I__803 (
            .O(N__4176),
            .I(N__4149));
    LocalMux I__802 (
            .O(N__4173),
            .I(N__4146));
    InMux I__801 (
            .O(N__4172),
            .I(N__4141));
    InMux I__800 (
            .O(N__4169),
            .I(N__4141));
    LocalMux I__799 (
            .O(N__4166),
            .I(N__4132));
    LocalMux I__798 (
            .O(N__4161),
            .I(N__4132));
    Span4Mux_h I__797 (
            .O(N__4158),
            .I(N__4132));
    LocalMux I__796 (
            .O(N__4155),
            .I(N__4132));
    Span4Mux_h I__795 (
            .O(N__4152),
            .I(N__4129));
    Odrv4 I__794 (
            .O(N__4149),
            .I(delayConstantZ0Z_2));
    Odrv12 I__793 (
            .O(N__4146),
            .I(delayConstantZ0Z_2));
    LocalMux I__792 (
            .O(N__4141),
            .I(delayConstantZ0Z_2));
    Odrv4 I__791 (
            .O(N__4132),
            .I(delayConstantZ0Z_2));
    Odrv4 I__790 (
            .O(N__4129),
            .I(delayConstantZ0Z_2));
    CascadeMux I__789 (
            .O(N__4118),
            .I(\dig1.m47_ns_1_cascade_ ));
    InMux I__788 (
            .O(N__4115),
            .I(N__4108));
    InMux I__787 (
            .O(N__4114),
            .I(N__4105));
    InMux I__786 (
            .O(N__4113),
            .I(N__4102));
    InMux I__785 (
            .O(N__4112),
            .I(N__4099));
    InMux I__784 (
            .O(N__4111),
            .I(N__4096));
    LocalMux I__783 (
            .O(N__4108),
            .I(N__4093));
    LocalMux I__782 (
            .O(N__4105),
            .I(col_1_1));
    LocalMux I__781 (
            .O(N__4102),
            .I(col_1_1));
    LocalMux I__780 (
            .O(N__4099),
            .I(col_1_1));
    LocalMux I__779 (
            .O(N__4096),
            .I(col_1_1));
    Odrv4 I__778 (
            .O(N__4093),
            .I(col_1_1));
    InMux I__777 (
            .O(N__4082),
            .I(N__4079));
    LocalMux I__776 (
            .O(N__4079),
            .I(\dig1.N_49 ));
    InMux I__775 (
            .O(N__4076),
            .I(N__4073));
    LocalMux I__774 (
            .O(N__4073),
            .I(\dig1.m41_bm ));
    CascadeMux I__773 (
            .O(N__4070),
            .I(\dig1.m41_am_cascade_ ));
    InMux I__772 (
            .O(N__4067),
            .I(N__4064));
    LocalMux I__771 (
            .O(N__4064),
            .I(\dig1.N_44 ));
    CascadeMux I__770 (
            .O(N__4061),
            .I(\dig1.m10_ns_1_cascade_ ));
    InMux I__769 (
            .O(N__4058),
            .I(N__4055));
    LocalMux I__768 (
            .O(N__4055),
            .I(\dig1.N_11_0 ));
    InMux I__767 (
            .O(N__4052),
            .I(N__4041));
    InMux I__766 (
            .O(N__4051),
            .I(N__4041));
    CascadeMux I__765 (
            .O(N__4050),
            .I(N__4033));
    InMux I__764 (
            .O(N__4049),
            .I(N__4028));
    InMux I__763 (
            .O(N__4048),
            .I(N__4028));
    InMux I__762 (
            .O(N__4047),
            .I(N__4023));
    InMux I__761 (
            .O(N__4046),
            .I(N__4023));
    LocalMux I__760 (
            .O(N__4041),
            .I(N__4020));
    InMux I__759 (
            .O(N__4040),
            .I(N__4015));
    InMux I__758 (
            .O(N__4039),
            .I(N__4015));
    InMux I__757 (
            .O(N__4038),
            .I(N__4010));
    InMux I__756 (
            .O(N__4037),
            .I(N__4010));
    InMux I__755 (
            .O(N__4036),
            .I(N__4007));
    InMux I__754 (
            .O(N__4033),
            .I(N__4004));
    LocalMux I__753 (
            .O(N__4028),
            .I(N__3999));
    LocalMux I__752 (
            .O(N__4023),
            .I(N__3999));
    Sp12to4 I__751 (
            .O(N__4020),
            .I(N__3992));
    LocalMux I__750 (
            .O(N__4015),
            .I(N__3992));
    LocalMux I__749 (
            .O(N__4010),
            .I(N__3992));
    LocalMux I__748 (
            .O(N__4007),
            .I(delayConstantZ0Z_6));
    LocalMux I__747 (
            .O(N__4004),
            .I(delayConstantZ0Z_6));
    Odrv4 I__746 (
            .O(N__3999),
            .I(delayConstantZ0Z_6));
    Odrv12 I__745 (
            .O(N__3992),
            .I(delayConstantZ0Z_6));
    InMux I__744 (
            .O(N__3983),
            .I(N__3980));
    LocalMux I__743 (
            .O(N__3980),
            .I(olddn_RNIM5BH1Z0Z_1));
    InMux I__742 (
            .O(N__3977),
            .I(un1_delayConstant_cry_0));
    InMux I__741 (
            .O(N__3974),
            .I(N__3971));
    LocalMux I__740 (
            .O(N__3971),
            .I(olddn_RNIM5BHZ0Z1));
    InMux I__739 (
            .O(N__3968),
            .I(un1_delayConstant_cry_1));
    CascadeMux I__738 (
            .O(N__3965),
            .I(N__3962));
    InMux I__737 (
            .O(N__3962),
            .I(N__3959));
    LocalMux I__736 (
            .O(N__3959),
            .I(olddn_RNIM5BH1Z0Z_2));
    InMux I__735 (
            .O(N__3956),
            .I(un1_delayConstant_cry_2));
    CascadeMux I__734 (
            .O(N__3953),
            .I(N__3950));
    InMux I__733 (
            .O(N__3950),
            .I(N__3947));
    LocalMux I__732 (
            .O(N__3947),
            .I(N__3944));
    Odrv4 I__731 (
            .O(N__3944),
            .I(olddn_RNIM5BH1Z0Z_3));
    InMux I__730 (
            .O(N__3941),
            .I(un1_delayConstant_cry_3));
    InMux I__729 (
            .O(N__3938),
            .I(N__3935));
    LocalMux I__728 (
            .O(N__3935),
            .I(olddn_RNIM5BH1Z0Z_0));
    InMux I__727 (
            .O(N__3932),
            .I(un1_delayConstant_cry_4));
    CascadeMux I__726 (
            .O(N__3929),
            .I(N__3926));
    InMux I__725 (
            .O(N__3926),
            .I(N__3923));
    LocalMux I__724 (
            .O(N__3923),
            .I(N__3920));
    Odrv4 I__723 (
            .O(N__3920),
            .I(olddn_RNIM5BH1Z0Z_4));
    InMux I__722 (
            .O(N__3917),
            .I(un1_delayConstant_cry_5));
    CascadeMux I__721 (
            .O(N__3914),
            .I(N__3908));
    InMux I__720 (
            .O(N__3913),
            .I(N__3901));
    InMux I__719 (
            .O(N__3912),
            .I(N__3898));
    InMux I__718 (
            .O(N__3911),
            .I(N__3891));
    InMux I__717 (
            .O(N__3908),
            .I(N__3891));
    InMux I__716 (
            .O(N__3907),
            .I(N__3891));
    InMux I__715 (
            .O(N__3906),
            .I(N__3884));
    InMux I__714 (
            .O(N__3905),
            .I(N__3884));
    InMux I__713 (
            .O(N__3904),
            .I(N__3884));
    LocalMux I__712 (
            .O(N__3901),
            .I(delayConstant16_i));
    LocalMux I__711 (
            .O(N__3898),
            .I(delayConstant16_i));
    LocalMux I__710 (
            .O(N__3891),
            .I(delayConstant16_i));
    LocalMux I__709 (
            .O(N__3884),
            .I(delayConstant16_i));
    InMux I__708 (
            .O(N__3875),
            .I(N__3864));
    InMux I__707 (
            .O(N__3874),
            .I(N__3861));
    InMux I__706 (
            .O(N__3873),
            .I(N__3854));
    InMux I__705 (
            .O(N__3872),
            .I(N__3854));
    InMux I__704 (
            .O(N__3871),
            .I(N__3854));
    InMux I__703 (
            .O(N__3870),
            .I(N__3845));
    InMux I__702 (
            .O(N__3869),
            .I(N__3845));
    InMux I__701 (
            .O(N__3868),
            .I(N__3845));
    InMux I__700 (
            .O(N__3867),
            .I(N__3845));
    LocalMux I__699 (
            .O(N__3864),
            .I(olddn_RNIEENHZ0));
    LocalMux I__698 (
            .O(N__3861),
            .I(olddn_RNIEENHZ0));
    LocalMux I__697 (
            .O(N__3854),
            .I(olddn_RNIEENHZ0));
    LocalMux I__696 (
            .O(N__3845),
            .I(olddn_RNIEENHZ0));
    InMux I__695 (
            .O(N__3836),
            .I(un1_delayConstant_cry_6));
    CascadeMux I__694 (
            .O(N__3833),
            .I(\dig1.N_15_cascade_ ));
    InMux I__693 (
            .O(N__3830),
            .I(N__3827));
    LocalMux I__692 (
            .O(N__3827),
            .I(\dig1.N_18 ));
    CascadeMux I__691 (
            .O(N__3824),
            .I(N__3821));
    InMux I__690 (
            .O(N__3821),
            .I(N__3816));
    InMux I__689 (
            .O(N__3820),
            .I(N__3813));
    InMux I__688 (
            .O(N__3819),
            .I(N__3808));
    LocalMux I__687 (
            .O(N__3816),
            .I(N__3803));
    LocalMux I__686 (
            .O(N__3813),
            .I(N__3803));
    InMux I__685 (
            .O(N__3812),
            .I(N__3800));
    InMux I__684 (
            .O(N__3811),
            .I(N__3797));
    LocalMux I__683 (
            .O(N__3808),
            .I(slowclk));
    Odrv4 I__682 (
            .O(N__3803),
            .I(slowclk));
    LocalMux I__681 (
            .O(N__3800),
            .I(slowclk));
    LocalMux I__680 (
            .O(N__3797),
            .I(slowclk));
    InMux I__679 (
            .O(N__3788),
            .I(N__3782));
    InMux I__678 (
            .O(N__3787),
            .I(N__3782));
    LocalMux I__677 (
            .O(N__3782),
            .I(clock_out_RNIR6ER));
    InMux I__676 (
            .O(N__3779),
            .I(N__3776));
    LocalMux I__675 (
            .O(N__3776),
            .I(\dig1.N_17 ));
    InMux I__674 (
            .O(N__3773),
            .I(N__3770));
    LocalMux I__673 (
            .O(N__3770),
            .I(\dig1.m32_bm ));
    CascadeMux I__672 (
            .O(N__3767),
            .I(N__3764));
    InMux I__671 (
            .O(N__3764),
            .I(N__3761));
    LocalMux I__670 (
            .O(N__3761),
            .I(\dig1.m32_am ));
    IoInMux I__669 (
            .O(N__3758),
            .I(N__3755));
    LocalMux I__668 (
            .O(N__3755),
            .I(N__3752));
    Span4Mux_s2_v I__667 (
            .O(N__3752),
            .I(N__3749));
    Sp12to4 I__666 (
            .O(N__3749),
            .I(N__3746));
    Span12Mux_h I__665 (
            .O(N__3746),
            .I(N__3743));
    Span12Mux_v I__664 (
            .O(N__3743),
            .I(N__3740));
    Odrv12 I__663 (
            .O(N__3740),
            .I(leds_1_i_2));
    CascadeMux I__662 (
            .O(N__3737),
            .I(N__3734));
    InMux I__661 (
            .O(N__3734),
            .I(N__3731));
    LocalMux I__660 (
            .O(N__3731),
            .I(un1_delayConstant_cry_0_c_RNOZ0));
    InMux I__659 (
            .O(N__3728),
            .I(N__3725));
    LocalMux I__658 (
            .O(N__3725),
            .I(\dig1.m77_am ));
    InMux I__657 (
            .O(N__3722),
            .I(N__3719));
    LocalMux I__656 (
            .O(N__3719),
            .I(N__3716));
    Span4Mux_h I__655 (
            .O(N__3716),
            .I(N__3713));
    Odrv4 I__654 (
            .O(N__3713),
            .I(\debounceup.out_cnv_2 ));
    CascadeMux I__653 (
            .O(N__3710),
            .I(N__3707));
    InMux I__652 (
            .O(N__3707),
            .I(N__3704));
    LocalMux I__651 (
            .O(N__3704),
            .I(N__3701));
    Span12Mux_h I__650 (
            .O(N__3701),
            .I(N__3698));
    Span12Mux_v I__649 (
            .O(N__3698),
            .I(N__3695));
    Odrv12 I__648 (
            .O(N__3695),
            .I(delup_c));
    InMux I__647 (
            .O(N__3692),
            .I(N__3687));
    InMux I__646 (
            .O(N__3691),
            .I(N__3682));
    InMux I__645 (
            .O(N__3690),
            .I(N__3682));
    LocalMux I__644 (
            .O(N__3687),
            .I(debouncedup));
    LocalMux I__643 (
            .O(N__3682),
            .I(debouncedup));
    InMux I__642 (
            .O(N__3677),
            .I(N__3674));
    LocalMux I__641 (
            .O(N__3674),
            .I(N__3671));
    Odrv4 I__640 (
            .O(N__3671),
            .I(\dig1.m77_bm ));
    IoInMux I__639 (
            .O(N__3668),
            .I(N__3665));
    LocalMux I__638 (
            .O(N__3665),
            .I(N__3662));
    IoSpan4Mux I__637 (
            .O(N__3662),
            .I(N__3659));
    IoSpan4Mux I__636 (
            .O(N__3659),
            .I(N__3656));
    Sp12to4 I__635 (
            .O(N__3656),
            .I(N__3653));
    Span12Mux_s6_v I__634 (
            .O(N__3653),
            .I(N__3650));
    Odrv12 I__633 (
            .O(N__3650),
            .I(leds_1_i_1));
    IoInMux I__632 (
            .O(N__3647),
            .I(N__3644));
    LocalMux I__631 (
            .O(N__3644),
            .I(N__3641));
    Span12Mux_s5_v I__630 (
            .O(N__3641),
            .I(N__3638));
    Span12Mux_v I__629 (
            .O(N__3638),
            .I(N__3635));
    Odrv12 I__628 (
            .O(N__3635),
            .I(lcol1_c));
    InMux I__627 (
            .O(N__3632),
            .I(N__3629));
    LocalMux I__626 (
            .O(N__3629),
            .I(\dig1.N_39 ));
    IoInMux I__625 (
            .O(N__3626),
            .I(N__3623));
    LocalMux I__624 (
            .O(N__3623),
            .I(N__3620));
    IoSpan4Mux I__623 (
            .O(N__3620),
            .I(N__3617));
    Span4Mux_s3_v I__622 (
            .O(N__3617),
            .I(N__3614));
    Sp12to4 I__621 (
            .O(N__3614),
            .I(N__3611));
    Span12Mux_s10_v I__620 (
            .O(N__3611),
            .I(N__3608));
    Span12Mux_h I__619 (
            .O(N__3608),
            .I(N__3605));
    Odrv12 I__618 (
            .O(N__3605),
            .I(leds_1_i_3));
    IoInMux I__617 (
            .O(N__3602),
            .I(N__3599));
    LocalMux I__616 (
            .O(N__3599),
            .I(N__3596));
    IoSpan4Mux I__615 (
            .O(N__3596),
            .I(N__3592));
    InMux I__614 (
            .O(N__3595),
            .I(N__3589));
    Span4Mux_s2_v I__613 (
            .O(N__3592),
            .I(N__3586));
    LocalMux I__612 (
            .O(N__3589),
            .I(N__3580));
    Span4Mux_v I__611 (
            .O(N__3586),
            .I(N__3577));
    InMux I__610 (
            .O(N__3585),
            .I(N__3574));
    InMux I__609 (
            .O(N__3584),
            .I(N__3571));
    InMux I__608 (
            .O(N__3583),
            .I(N__3568));
    Span4Mux_v I__607 (
            .O(N__3580),
            .I(N__3565));
    Span4Mux_v I__606 (
            .O(N__3577),
            .I(N__3560));
    LocalMux I__605 (
            .O(N__3574),
            .I(N__3560));
    LocalMux I__604 (
            .O(N__3571),
            .I(N__3554));
    LocalMux I__603 (
            .O(N__3568),
            .I(N__3554));
    Span4Mux_h I__602 (
            .O(N__3565),
            .I(N__3549));
    Span4Mux_v I__601 (
            .O(N__3560),
            .I(N__3549));
    InMux I__600 (
            .O(N__3559),
            .I(N__3546));
    Span4Mux_v I__599 (
            .O(N__3554),
            .I(N__3543));
    Sp12to4 I__598 (
            .O(N__3549),
            .I(N__3538));
    LocalMux I__597 (
            .O(N__3546),
            .I(N__3538));
    Sp12to4 I__596 (
            .O(N__3543),
            .I(N__3535));
    Span12Mux_h I__595 (
            .O(N__3538),
            .I(N__3532));
    Span12Mux_h I__594 (
            .O(N__3535),
            .I(N__3529));
    Span12Mux_v I__593 (
            .O(N__3532),
            .I(N__3526));
    Span12Mux_v I__592 (
            .O(N__3529),
            .I(N__3523));
    Odrv12 I__591 (
            .O(N__3526),
            .I(masterreset_c));
    Odrv12 I__590 (
            .O(N__3523),
            .I(masterreset_c));
    CascadeMux I__589 (
            .O(N__3518),
            .I(delayConstant16_i_cascade_));
    InMux I__588 (
            .O(N__3515),
            .I(N__3512));
    LocalMux I__587 (
            .O(N__3512),
            .I(oldupZ0));
    CascadeMux I__586 (
            .O(N__3509),
            .I(N__3506));
    InMux I__585 (
            .O(N__3506),
            .I(N__3501));
    InMux I__584 (
            .O(N__3505),
            .I(N__3496));
    InMux I__583 (
            .O(N__3504),
            .I(N__3496));
    LocalMux I__582 (
            .O(N__3501),
            .I(debounceddn));
    LocalMux I__581 (
            .O(N__3496),
            .I(debounceddn));
    InMux I__580 (
            .O(N__3491),
            .I(N__3488));
    LocalMux I__579 (
            .O(N__3488),
            .I(olddnZ0));
    InMux I__578 (
            .O(N__3485),
            .I(N__3482));
    LocalMux I__577 (
            .O(N__3482),
            .I(\dig1.N_72 ));
    InMux I__576 (
            .O(N__3479),
            .I(N__3476));
    LocalMux I__575 (
            .O(N__3476),
            .I(N__3473));
    Span4Mux_h I__574 (
            .O(N__3473),
            .I(N__3470));
    Odrv4 I__573 (
            .O(N__3470),
            .I(\debouncedn.out_cnv_2 ));
    InMux I__572 (
            .O(N__3467),
            .I(N__3464));
    LocalMux I__571 (
            .O(N__3464),
            .I(N__3461));
    Span4Mux_v I__570 (
            .O(N__3461),
            .I(N__3458));
    Sp12to4 I__569 (
            .O(N__3458),
            .I(N__3455));
    Span12Mux_h I__568 (
            .O(N__3455),
            .I(N__3452));
    Span12Mux_v I__567 (
            .O(N__3452),
            .I(N__3449));
    Odrv12 I__566 (
            .O(N__3449),
            .I(deldn_c));
    CascadeMux I__565 (
            .O(N__3446),
            .I(\dig1.N_58_cascade_ ));
    InMux I__564 (
            .O(N__3443),
            .I(N__3440));
    LocalMux I__563 (
            .O(N__3440),
            .I(\dig1.leds_17_i_ns_1_2 ));
    InMux I__562 (
            .O(N__3437),
            .I(N__3434));
    LocalMux I__561 (
            .O(N__3434),
            .I(\dig1.N_61 ));
    InMux I__560 (
            .O(N__3431),
            .I(N__3428));
    LocalMux I__559 (
            .O(N__3428),
            .I(\dig1.m68_bm ));
    InMux I__558 (
            .O(N__3425),
            .I(N__3422));
    LocalMux I__557 (
            .O(N__3422),
            .I(\dig1.m68_am ));
    InMux I__556 (
            .O(N__3419),
            .I(N__3402));
    InMux I__555 (
            .O(N__3418),
            .I(N__3399));
    InMux I__554 (
            .O(N__3417),
            .I(N__3390));
    InMux I__553 (
            .O(N__3416),
            .I(N__3390));
    InMux I__552 (
            .O(N__3415),
            .I(N__3390));
    InMux I__551 (
            .O(N__3414),
            .I(N__3381));
    InMux I__550 (
            .O(N__3413),
            .I(N__3381));
    InMux I__549 (
            .O(N__3412),
            .I(N__3381));
    InMux I__548 (
            .O(N__3411),
            .I(N__3381));
    InMux I__547 (
            .O(N__3410),
            .I(N__3374));
    InMux I__546 (
            .O(N__3409),
            .I(N__3374));
    InMux I__545 (
            .O(N__3408),
            .I(N__3374));
    InMux I__544 (
            .O(N__3407),
            .I(N__3367));
    InMux I__543 (
            .O(N__3406),
            .I(N__3367));
    InMux I__542 (
            .O(N__3405),
            .I(N__3367));
    LocalMux I__541 (
            .O(N__3402),
            .I(N__3362));
    LocalMux I__540 (
            .O(N__3399),
            .I(N__3362));
    InMux I__539 (
            .O(N__3398),
            .I(N__3359));
    InMux I__538 (
            .O(N__3397),
            .I(N__3356));
    LocalMux I__537 (
            .O(N__3390),
            .I(\arses.counter8 ));
    LocalMux I__536 (
            .O(N__3381),
            .I(\arses.counter8 ));
    LocalMux I__535 (
            .O(N__3374),
            .I(\arses.counter8 ));
    LocalMux I__534 (
            .O(N__3367),
            .I(\arses.counter8 ));
    Odrv4 I__533 (
            .O(N__3362),
            .I(\arses.counter8 ));
    LocalMux I__532 (
            .O(N__3359),
            .I(\arses.counter8 ));
    LocalMux I__531 (
            .O(N__3356),
            .I(\arses.counter8 ));
    IoInMux I__530 (
            .O(N__3341),
            .I(N__3338));
    LocalMux I__529 (
            .O(N__3338),
            .I(N__3335));
    IoSpan4Mux I__528 (
            .O(N__3335),
            .I(N__3332));
    Span4Mux_s3_v I__527 (
            .O(N__3332),
            .I(N__3329));
    Sp12to4 I__526 (
            .O(N__3329),
            .I(N__3326));
    Span12Mux_h I__525 (
            .O(N__3326),
            .I(N__3323));
    Span12Mux_v I__524 (
            .O(N__3323),
            .I(N__3320));
    Odrv12 I__523 (
            .O(N__3320),
            .I(lcol2_c));
    InMux I__522 (
            .O(N__3317),
            .I(N__3313));
    InMux I__521 (
            .O(N__3316),
            .I(N__3310));
    LocalMux I__520 (
            .O(N__3313),
            .I(\arses.counterZ0Z_7 ));
    LocalMux I__519 (
            .O(N__3310),
            .I(\arses.counterZ0Z_7 ));
    InMux I__518 (
            .O(N__3305),
            .I(N__3301));
    InMux I__517 (
            .O(N__3304),
            .I(N__3298));
    LocalMux I__516 (
            .O(N__3301),
            .I(\arses.counterZ0Z_6 ));
    LocalMux I__515 (
            .O(N__3298),
            .I(\arses.counterZ0Z_6 ));
    CascadeMux I__514 (
            .O(N__3293),
            .I(N__3289));
    InMux I__513 (
            .O(N__3292),
            .I(N__3286));
    InMux I__512 (
            .O(N__3289),
            .I(N__3283));
    LocalMux I__511 (
            .O(N__3286),
            .I(\arses.counterZ0Z_8 ));
    LocalMux I__510 (
            .O(N__3283),
            .I(\arses.counterZ0Z_8 ));
    InMux I__509 (
            .O(N__3278),
            .I(N__3274));
    InMux I__508 (
            .O(N__3277),
            .I(N__3271));
    LocalMux I__507 (
            .O(N__3274),
            .I(\arses.counterZ0Z_5 ));
    LocalMux I__506 (
            .O(N__3271),
            .I(\arses.counterZ0Z_5 ));
    InMux I__505 (
            .O(N__3266),
            .I(N__3262));
    InMux I__504 (
            .O(N__3265),
            .I(N__3259));
    LocalMux I__503 (
            .O(N__3262),
            .I(\arses.counterZ0Z_4 ));
    LocalMux I__502 (
            .O(N__3259),
            .I(\arses.counterZ0Z_4 ));
    InMux I__501 (
            .O(N__3254),
            .I(N__3249));
    InMux I__500 (
            .O(N__3253),
            .I(N__3246));
    InMux I__499 (
            .O(N__3252),
            .I(N__3243));
    LocalMux I__498 (
            .O(N__3249),
            .I(N__3240));
    LocalMux I__497 (
            .O(N__3246),
            .I(N__3237));
    LocalMux I__496 (
            .O(N__3243),
            .I(\arses.counterZ0Z_1 ));
    Odrv4 I__495 (
            .O(N__3240),
            .I(\arses.counterZ0Z_1 ));
    Odrv4 I__494 (
            .O(N__3237),
            .I(\arses.counterZ0Z_1 ));
    CascadeMux I__493 (
            .O(N__3230),
            .I(\arses.un1_counterlto8_2_cascade_ ));
    InMux I__492 (
            .O(N__3227),
            .I(N__3223));
    InMux I__491 (
            .O(N__3226),
            .I(N__3220));
    LocalMux I__490 (
            .O(N__3223),
            .I(\arses.counterZ0Z_11 ));
    LocalMux I__489 (
            .O(N__3220),
            .I(\arses.counterZ0Z_11 ));
    InMux I__488 (
            .O(N__3215),
            .I(N__3211));
    InMux I__487 (
            .O(N__3214),
            .I(N__3208));
    LocalMux I__486 (
            .O(N__3211),
            .I(\arses.counterZ0Z_10 ));
    LocalMux I__485 (
            .O(N__3208),
            .I(\arses.counterZ0Z_10 ));
    CascadeMux I__484 (
            .O(N__3203),
            .I(\arses.un1_counterlt11_cascade_ ));
    InMux I__483 (
            .O(N__3200),
            .I(N__3196));
    InMux I__482 (
            .O(N__3199),
            .I(N__3193));
    LocalMux I__481 (
            .O(N__3196),
            .I(\arses.counterZ0Z_9 ));
    LocalMux I__480 (
            .O(N__3193),
            .I(\arses.counterZ0Z_9 ));
    InMux I__479 (
            .O(N__3188),
            .I(N__3184));
    InMux I__478 (
            .O(N__3187),
            .I(N__3181));
    LocalMux I__477 (
            .O(N__3184),
            .I(\arses.counterZ0Z_14 ));
    LocalMux I__476 (
            .O(N__3181),
            .I(\arses.counterZ0Z_14 ));
    InMux I__475 (
            .O(N__3176),
            .I(N__3172));
    InMux I__474 (
            .O(N__3175),
            .I(N__3169));
    LocalMux I__473 (
            .O(N__3172),
            .I(\arses.counterZ0Z_13 ));
    LocalMux I__472 (
            .O(N__3169),
            .I(\arses.counterZ0Z_13 ));
    CascadeMux I__471 (
            .O(N__3164),
            .I(\arses.un1_counterlt13_0_cascade_ ));
    InMux I__470 (
            .O(N__3161),
            .I(N__3157));
    InMux I__469 (
            .O(N__3160),
            .I(N__3154));
    LocalMux I__468 (
            .O(N__3157),
            .I(\arses.counterZ0Z_12 ));
    LocalMux I__467 (
            .O(N__3154),
            .I(\arses.counterZ0Z_12 ));
    CascadeMux I__466 (
            .O(N__3149),
            .I(\arses.counter8_cascade_ ));
    InMux I__465 (
            .O(N__3146),
            .I(N__3142));
    InMux I__464 (
            .O(N__3145),
            .I(N__3139));
    LocalMux I__463 (
            .O(N__3142),
            .I(\arses.counterZ0Z_3 ));
    LocalMux I__462 (
            .O(N__3139),
            .I(\arses.counterZ0Z_3 ));
    InMux I__461 (
            .O(N__3134),
            .I(N__3130));
    InMux I__460 (
            .O(N__3133),
            .I(N__3127));
    LocalMux I__459 (
            .O(N__3130),
            .I(\arses.counterZ0Z_2 ));
    LocalMux I__458 (
            .O(N__3127),
            .I(\arses.counterZ0Z_2 ));
    InMux I__457 (
            .O(N__3122),
            .I(N__3119));
    LocalMux I__456 (
            .O(N__3119),
            .I(\arses.un1_counterlto4_2 ));
    CascadeMux I__455 (
            .O(N__3116),
            .I(N__3113));
    InMux I__454 (
            .O(N__3113),
            .I(N__3108));
    InMux I__453 (
            .O(N__3112),
            .I(N__3104));
    InMux I__452 (
            .O(N__3111),
            .I(N__3101));
    LocalMux I__451 (
            .O(N__3108),
            .I(N__3098));
    InMux I__450 (
            .O(N__3107),
            .I(N__3095));
    LocalMux I__449 (
            .O(N__3104),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__448 (
            .O(N__3101),
            .I(\arses.counterZ0Z_0 ));
    Odrv4 I__447 (
            .O(N__3098),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__446 (
            .O(N__3095),
            .I(\arses.counterZ0Z_0 ));
    InMux I__445 (
            .O(N__3086),
            .I(N__3083));
    LocalMux I__444 (
            .O(N__3083),
            .I(\dig1.N_78 ));
    InMux I__443 (
            .O(N__3080),
            .I(\arses.un2_counter_cry_13 ));
    IoInMux I__442 (
            .O(N__3077),
            .I(N__3074));
    LocalMux I__441 (
            .O(N__3074),
            .I(N__3071));
    IoSpan4Mux I__440 (
            .O(N__3071),
            .I(N__3068));
    IoSpan4Mux I__439 (
            .O(N__3068),
            .I(N__3065));
    Span4Mux_s3_v I__438 (
            .O(N__3065),
            .I(N__3062));
    Sp12to4 I__437 (
            .O(N__3062),
            .I(N__3059));
    Span12Mux_s11_v I__436 (
            .O(N__3059),
            .I(N__3056));
    Odrv12 I__435 (
            .O(N__3056),
            .I(leds_1_i_0_3));
    CascadeMux I__434 (
            .O(N__3053),
            .I(\debounceup.counter_RNI45V02Z0Z_4_cascade_ ));
    InMux I__433 (
            .O(N__3050),
            .I(N__3042));
    InMux I__432 (
            .O(N__3049),
            .I(N__3042));
    InMux I__431 (
            .O(N__3048),
            .I(N__3039));
    InMux I__430 (
            .O(N__3047),
            .I(N__3036));
    LocalMux I__429 (
            .O(N__3042),
            .I(\debounceup.counterZ0Z_3 ));
    LocalMux I__428 (
            .O(N__3039),
            .I(\debounceup.counterZ0Z_3 ));
    LocalMux I__427 (
            .O(N__3036),
            .I(\debounceup.counterZ0Z_3 ));
    InMux I__426 (
            .O(N__3029),
            .I(N__3021));
    InMux I__425 (
            .O(N__3028),
            .I(N__3021));
    InMux I__424 (
            .O(N__3027),
            .I(N__3016));
    InMux I__423 (
            .O(N__3026),
            .I(N__3016));
    LocalMux I__422 (
            .O(N__3021),
            .I(\debounceup.counterZ0Z_2 ));
    LocalMux I__421 (
            .O(N__3016),
            .I(\debounceup.counterZ0Z_2 ));
    InMux I__420 (
            .O(N__3011),
            .I(N__3006));
    InMux I__419 (
            .O(N__3010),
            .I(N__3001));
    InMux I__418 (
            .O(N__3009),
            .I(N__3001));
    LocalMux I__417 (
            .O(N__3006),
            .I(\debounceup.counterZ0Z_4 ));
    LocalMux I__416 (
            .O(N__3001),
            .I(\debounceup.counterZ0Z_4 ));
    CascadeMux I__415 (
            .O(N__2996),
            .I(\debounceup.counter18_0_2_cascade_ ));
    CascadeMux I__414 (
            .O(N__2993),
            .I(N__2989));
    CascadeMux I__413 (
            .O(N__2992),
            .I(N__2985));
    InMux I__412 (
            .O(N__2989),
            .I(N__2981));
    InMux I__411 (
            .O(N__2988),
            .I(N__2974));
    InMux I__410 (
            .O(N__2985),
            .I(N__2974));
    InMux I__409 (
            .O(N__2984),
            .I(N__2974));
    LocalMux I__408 (
            .O(N__2981),
            .I(\debounceup.counterZ0Z_0 ));
    LocalMux I__407 (
            .O(N__2974),
            .I(\debounceup.counterZ0Z_0 ));
    CascadeMux I__406 (
            .O(N__2969),
            .I(N__2966));
    InMux I__405 (
            .O(N__2966),
            .I(N__2962));
    InMux I__404 (
            .O(N__2965),
            .I(N__2957));
    LocalMux I__403 (
            .O(N__2962),
            .I(N__2954));
    InMux I__402 (
            .O(N__2961),
            .I(N__2949));
    InMux I__401 (
            .O(N__2960),
            .I(N__2949));
    LocalMux I__400 (
            .O(N__2957),
            .I(\debounceup.counter_RNI45V02Z0Z_4 ));
    Odrv4 I__399 (
            .O(N__2954),
            .I(\debounceup.counter_RNI45V02Z0Z_4 ));
    LocalMux I__398 (
            .O(N__2949),
            .I(\debounceup.counter_RNI45V02Z0Z_4 ));
    InMux I__397 (
            .O(N__2942),
            .I(N__2935));
    InMux I__396 (
            .O(N__2941),
            .I(N__2935));
    InMux I__395 (
            .O(N__2940),
            .I(N__2932));
    LocalMux I__394 (
            .O(N__2935),
            .I(\debounceup.counterZ0Z_1 ));
    LocalMux I__393 (
            .O(N__2932),
            .I(\debounceup.counterZ0Z_1 ));
    IoInMux I__392 (
            .O(N__2927),
            .I(N__2924));
    LocalMux I__391 (
            .O(N__2924),
            .I(N__2921));
    IoSpan4Mux I__390 (
            .O(N__2921),
            .I(N__2918));
    Span4Mux_s3_v I__389 (
            .O(N__2918),
            .I(N__2915));
    Span4Mux_v I__388 (
            .O(N__2915),
            .I(N__2912));
    Sp12to4 I__387 (
            .O(N__2912),
            .I(N__2909));
    Span12Mux_v I__386 (
            .O(N__2909),
            .I(N__2906));
    Odrv12 I__385 (
            .O(N__2906),
            .I(leds_1_i_0_2));
    InMux I__384 (
            .O(N__2903),
            .I(\arses.un2_counter_cry_3 ));
    InMux I__383 (
            .O(N__2900),
            .I(\arses.un2_counter_cry_4 ));
    InMux I__382 (
            .O(N__2897),
            .I(\arses.un2_counter_cry_5 ));
    InMux I__381 (
            .O(N__2894),
            .I(\arses.un2_counter_cry_6 ));
    InMux I__380 (
            .O(N__2891),
            .I(\arses.un2_counter_cry_7 ));
    InMux I__379 (
            .O(N__2888),
            .I(bfn_17_17_0_));
    InMux I__378 (
            .O(N__2885),
            .I(\arses.un2_counter_cry_9 ));
    InMux I__377 (
            .O(N__2882),
            .I(\arses.un2_counter_cry_10 ));
    InMux I__376 (
            .O(N__2879),
            .I(\arses.un2_counter_cry_11 ));
    InMux I__375 (
            .O(N__2876),
            .I(\arses.un2_counter_cry_12 ));
    InMux I__374 (
            .O(N__2873),
            .I(\debounceconsolereset.un3_counter_cry_3 ));
    InMux I__373 (
            .O(N__2870),
            .I(N__2865));
    InMux I__372 (
            .O(N__2869),
            .I(N__2860));
    InMux I__371 (
            .O(N__2868),
            .I(N__2860));
    LocalMux I__370 (
            .O(N__2865),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    LocalMux I__369 (
            .O(N__2860),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    CascadeMux I__368 (
            .O(N__2855),
            .I(clock_out_RNIR6ER_0_cascade_));
    InMux I__367 (
            .O(N__2852),
            .I(N__2849));
    LocalMux I__366 (
            .O(N__2849),
            .I(\debounceconsolereset.un3_counter_cry_2_THRU_CO ));
    CascadeMux I__365 (
            .O(N__2846),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4_cascade_ ));
    CascadeMux I__364 (
            .O(N__2843),
            .I(N__2838));
    CascadeMux I__363 (
            .O(N__2842),
            .I(N__2834));
    InMux I__362 (
            .O(N__2841),
            .I(N__2831));
    InMux I__361 (
            .O(N__2838),
            .I(N__2826));
    InMux I__360 (
            .O(N__2837),
            .I(N__2826));
    InMux I__359 (
            .O(N__2834),
            .I(N__2823));
    LocalMux I__358 (
            .O(N__2831),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    LocalMux I__357 (
            .O(N__2826),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    LocalMux I__356 (
            .O(N__2823),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    CascadeMux I__355 (
            .O(N__2816),
            .I(N__2812));
    InMux I__354 (
            .O(N__2815),
            .I(N__2807));
    InMux I__353 (
            .O(N__2812),
            .I(N__2804));
    InMux I__352 (
            .O(N__2811),
            .I(N__2799));
    InMux I__351 (
            .O(N__2810),
            .I(N__2799));
    LocalMux I__350 (
            .O(N__2807),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4 ));
    LocalMux I__349 (
            .O(N__2804),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4 ));
    LocalMux I__348 (
            .O(N__2799),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4 ));
    CascadeMux I__347 (
            .O(N__2792),
            .I(N__2789));
    InMux I__346 (
            .O(N__2789),
            .I(N__2786));
    LocalMux I__345 (
            .O(N__2786),
            .I(\debounceconsolereset.un3_counter_cry_1_THRU_CO ));
    InMux I__344 (
            .O(N__2783),
            .I(N__2777));
    InMux I__343 (
            .O(N__2782),
            .I(N__2772));
    InMux I__342 (
            .O(N__2781),
            .I(N__2772));
    InMux I__341 (
            .O(N__2780),
            .I(N__2769));
    LocalMux I__340 (
            .O(N__2777),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    LocalMux I__339 (
            .O(N__2772),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    LocalMux I__338 (
            .O(N__2769),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    InMux I__337 (
            .O(N__2762),
            .I(\arses.un2_counter_cry_1 ));
    InMux I__336 (
            .O(N__2759),
            .I(\arses.un2_counter_cry_2 ));
    InMux I__335 (
            .O(N__2756),
            .I(\debounceup.un3_counter_cry_1 ));
    InMux I__334 (
            .O(N__2753),
            .I(\debounceup.un3_counter_cry_2 ));
    InMux I__333 (
            .O(N__2750),
            .I(\debounceup.un3_counter_cry_3 ));
    InMux I__332 (
            .O(N__2747),
            .I(N__2744));
    LocalMux I__331 (
            .O(N__2744),
            .I(\debounceup.un3_counter_cry_2_THRU_CO ));
    InMux I__330 (
            .O(N__2741),
            .I(N__2738));
    LocalMux I__329 (
            .O(N__2738),
            .I(\debounceup.un3_counter_cry_1_THRU_CO ));
    InMux I__328 (
            .O(N__2735),
            .I(N__2728));
    InMux I__327 (
            .O(N__2734),
            .I(N__2728));
    InMux I__326 (
            .O(N__2733),
            .I(N__2725));
    LocalMux I__325 (
            .O(N__2728),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    LocalMux I__324 (
            .O(N__2725),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    CascadeMux I__323 (
            .O(N__2720),
            .I(N__2716));
    CascadeMux I__322 (
            .O(N__2719),
            .I(N__2711));
    InMux I__321 (
            .O(N__2716),
            .I(N__2704));
    InMux I__320 (
            .O(N__2715),
            .I(N__2704));
    InMux I__319 (
            .O(N__2714),
            .I(N__2704));
    InMux I__318 (
            .O(N__2711),
            .I(N__2701));
    LocalMux I__317 (
            .O(N__2704),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    LocalMux I__316 (
            .O(N__2701),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    InMux I__315 (
            .O(N__2696),
            .I(\debounceconsolereset.un3_counter_cry_1 ));
    InMux I__314 (
            .O(N__2693),
            .I(\debounceconsolereset.un3_counter_cry_2 ));
    CascadeMux I__313 (
            .O(N__2690),
            .I(\debouncedn.counter_RNIBTPA2Z0Z_4_cascade_ ));
    CascadeMux I__312 (
            .O(N__2687),
            .I(N__2681));
    InMux I__311 (
            .O(N__2686),
            .I(N__2678));
    InMux I__310 (
            .O(N__2685),
            .I(N__2673));
    InMux I__309 (
            .O(N__2684),
            .I(N__2673));
    InMux I__308 (
            .O(N__2681),
            .I(N__2670));
    LocalMux I__307 (
            .O(N__2678),
            .I(\debouncedn.counterZ0Z_0 ));
    LocalMux I__306 (
            .O(N__2673),
            .I(\debouncedn.counterZ0Z_0 ));
    LocalMux I__305 (
            .O(N__2670),
            .I(\debouncedn.counterZ0Z_0 ));
    CascadeMux I__304 (
            .O(N__2663),
            .I(\debounceconsolereset.counter18_0_2_cascade_ ));
    InMux I__303 (
            .O(N__2660),
            .I(N__2657));
    LocalMux I__302 (
            .O(N__2657),
            .I(\debouncedn.un3_counter_cry_2_THRU_CO ));
    InMux I__301 (
            .O(N__2654),
            .I(N__2648));
    InMux I__300 (
            .O(N__2653),
            .I(N__2643));
    InMux I__299 (
            .O(N__2652),
            .I(N__2643));
    InMux I__298 (
            .O(N__2651),
            .I(N__2640));
    LocalMux I__297 (
            .O(N__2648),
            .I(\debouncedn.counterZ0Z_3 ));
    LocalMux I__296 (
            .O(N__2643),
            .I(\debouncedn.counterZ0Z_3 ));
    LocalMux I__295 (
            .O(N__2640),
            .I(\debouncedn.counterZ0Z_3 ));
    InMux I__294 (
            .O(N__2633),
            .I(N__2630));
    LocalMux I__293 (
            .O(N__2630),
            .I(\debouncedn.un3_counter_cry_1_THRU_CO ));
    CascadeMux I__292 (
            .O(N__2627),
            .I(N__2623));
    InMux I__291 (
            .O(N__2626),
            .I(N__2618));
    InMux I__290 (
            .O(N__2623),
            .I(N__2615));
    InMux I__289 (
            .O(N__2622),
            .I(N__2610));
    InMux I__288 (
            .O(N__2621),
            .I(N__2610));
    LocalMux I__287 (
            .O(N__2618),
            .I(\debouncedn.counter_RNIBTPA2Z0Z_4 ));
    LocalMux I__286 (
            .O(N__2615),
            .I(\debouncedn.counter_RNIBTPA2Z0Z_4 ));
    LocalMux I__285 (
            .O(N__2610),
            .I(\debouncedn.counter_RNIBTPA2Z0Z_4 ));
    InMux I__284 (
            .O(N__2603),
            .I(N__2595));
    InMux I__283 (
            .O(N__2602),
            .I(N__2595));
    InMux I__282 (
            .O(N__2601),
            .I(N__2592));
    InMux I__281 (
            .O(N__2600),
            .I(N__2589));
    LocalMux I__280 (
            .O(N__2595),
            .I(\debouncedn.counterZ0Z_2 ));
    LocalMux I__279 (
            .O(N__2592),
            .I(\debouncedn.counterZ0Z_2 ));
    LocalMux I__278 (
            .O(N__2589),
            .I(\debouncedn.counterZ0Z_2 ));
    InMux I__277 (
            .O(N__2582),
            .I(N__2579));
    LocalMux I__276 (
            .O(N__2579),
            .I(N__2576));
    Span4Mux_v I__275 (
            .O(N__2576),
            .I(N__2573));
    Sp12to4 I__274 (
            .O(N__2573),
            .I(N__2570));
    Span12Mux_h I__273 (
            .O(N__2570),
            .I(N__2567));
    Span12Mux_v I__272 (
            .O(N__2567),
            .I(N__2564));
    Odrv12 I__271 (
            .O(N__2564),
            .I(consolereset_c));
    InMux I__270 (
            .O(N__2561),
            .I(N__2558));
    LocalMux I__269 (
            .O(N__2558),
            .I(\debounceconsolereset.out_cnv_2 ));
    IoInMux I__268 (
            .O(N__2555),
            .I(N__2552));
    LocalMux I__267 (
            .O(N__2552),
            .I(N__2549));
    Sp12to4 I__266 (
            .O(N__2549),
            .I(N__2546));
    Span12Mux_s6_v I__265 (
            .O(N__2546),
            .I(N__2543));
    Odrv12 I__264 (
            .O(N__2543),
            .I(lcol3_c));
    IoInMux I__263 (
            .O(N__2540),
            .I(N__2537));
    LocalMux I__262 (
            .O(N__2537),
            .I(N__2534));
    IoSpan4Mux I__261 (
            .O(N__2534),
            .I(N__2531));
    IoSpan4Mux I__260 (
            .O(N__2531),
            .I(N__2528));
    Span4Mux_s3_v I__259 (
            .O(N__2528),
            .I(N__2525));
    Sp12to4 I__258 (
            .O(N__2525),
            .I(N__2522));
    Odrv12 I__257 (
            .O(N__2522),
            .I(lcol4_c));
    InMux I__256 (
            .O(N__2519),
            .I(\debouncedn.un3_counter_cry_1 ));
    InMux I__255 (
            .O(N__2516),
            .I(\debouncedn.un3_counter_cry_2 ));
    InMux I__254 (
            .O(N__2513),
            .I(\debouncedn.un3_counter_cry_3 ));
    IoInMux I__253 (
            .O(N__2510),
            .I(N__2507));
    LocalMux I__252 (
            .O(N__2507),
            .I(N__2504));
    IoSpan4Mux I__251 (
            .O(N__2504),
            .I(N__2501));
    Odrv4 I__250 (
            .O(N__2501),
            .I(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO));
    CascadeMux I__249 (
            .O(N__2498),
            .I(\debouncedn.counter18_0_2_cascade_ ));
    InMux I__248 (
            .O(N__2495),
            .I(N__2490));
    InMux I__247 (
            .O(N__2494),
            .I(N__2487));
    InMux I__246 (
            .O(N__2493),
            .I(N__2484));
    LocalMux I__245 (
            .O(N__2490),
            .I(\debouncedn.counterZ0Z_1 ));
    LocalMux I__244 (
            .O(N__2487),
            .I(\debouncedn.counterZ0Z_1 ));
    LocalMux I__243 (
            .O(N__2484),
            .I(\debouncedn.counterZ0Z_1 ));
    CascadeMux I__242 (
            .O(N__2477),
            .I(N__2472));
    InMux I__241 (
            .O(N__2476),
            .I(N__2469));
    InMux I__240 (
            .O(N__2475),
            .I(N__2466));
    InMux I__239 (
            .O(N__2472),
            .I(N__2463));
    LocalMux I__238 (
            .O(N__2469),
            .I(\debouncedn.counterZ0Z_4 ));
    LocalMux I__237 (
            .O(N__2466),
            .I(\debouncedn.counterZ0Z_4 ));
    LocalMux I__236 (
            .O(N__2463),
            .I(\debouncedn.counterZ0Z_4 ));
    IoInMux I__235 (
            .O(N__2456),
            .I(N__2453));
    LocalMux I__234 (
            .O(N__2453),
            .I(N__2450));
    IoSpan4Mux I__233 (
            .O(N__2450),
            .I(N__2447));
    Span4Mux_s2_v I__232 (
            .O(N__2447),
            .I(N__2444));
    Sp12to4 I__231 (
            .O(N__2444),
            .I(N__2441));
    Span12Mux_s10_v I__230 (
            .O(N__2441),
            .I(N__2438));
    Span12Mux_v I__229 (
            .O(N__2438),
            .I(N__2435));
    Span12Mux_h I__228 (
            .O(N__2435),
            .I(N__2432));
    Odrv12 I__227 (
            .O(N__2432),
            .I(\arse.divseven.io_0_D_IN_0 ));
    IoInMux I__226 (
            .O(N__2429),
            .I(N__2426));
    LocalMux I__225 (
            .O(N__2426),
            .I(N__2423));
    Span12Mux_s4_h I__224 (
            .O(N__2423),
            .I(N__2420));
    Odrv12 I__223 (
            .O(N__2420),
            .I(masterreset_c_i));
    ClkMux I__222 (
            .O(N__2417),
            .I(N__2414));
    GlobalMux I__221 (
            .O(N__2414),
            .I(N__2411));
    gio2CtrlBuf I__220 (
            .O(N__2411),
            .I(\arse.un1_io_0_1_g ));
    IoInMux I__219 (
            .O(N__2408),
            .I(N__2405));
    LocalMux I__218 (
            .O(N__2405),
            .I(N__2402));
    Span4Mux_s1_v I__217 (
            .O(N__2402),
            .I(N__2399));
    Sp12to4 I__216 (
            .O(N__2399),
            .I(N__2396));
    Span12Mux_h I__215 (
            .O(N__2396),
            .I(N__2393));
    Span12Mux_v I__214 (
            .O(N__2393),
            .I(N__2390));
    Span12Mux_v I__213 (
            .O(N__2390),
            .I(N__2387));
    Odrv12 I__212 (
            .O(N__2387),
            .I(\top_pll_nrtthrth.PLLOUTCORE ));
    INV \INVarse.divseven.dout_0C  (
            .O(\INVarse.divseven.dout_0C_net ),
            .I(N__5906));
    INV \INVarse.apuresetoutregC  (
            .O(\INVarse.apuresetoutregC_net ),
            .I(N__5913));
    INV \INVarse.apusynclatchedC  (
            .O(\INVarse.apusynclatchedC_net ),
            .I(N__2417));
    INV \INVarse.diveight.dout_0C  (
            .O(\INVarse.diveight.dout_0C_net ),
            .I(N__5911));
    INV \INVarse.doingsevenC  (
            .O(\INVarse.doingsevenC_net ),
            .I(N__5903));
    INV \INVarse.cpuclkresetC  (
            .O(\INVarse.cpuclkresetC_net ),
            .I(N__5907));
    INV \INVarse.cpuresetoutregC  (
            .O(\INVarse.cpuresetoutregC_net ),
            .I(N__5902));
    INV \INVarse.cpuresetcount_0C  (
            .O(\INVarse.cpuresetcount_0C_net ),
            .I(N__5901));
    defparam IN_MUX_bfv_21_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_12_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\arses.un2_counter_cry_8 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_27_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_27_8_0_));
    ICE_GB \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5  (
            .USERSIGNALTOGLOBALBUFFER(N__2408),
            .GLOBALBUFFEROUTPUT(PLLOUTCORE_g));
    ICE_GB \arse.divseven.io_0_RNIIG08  (
            .USERSIGNALTOGLOBALBUFFER(N__2456),
            .GLOBALBUFFEROUTPUT(\arse.un1_io_0_1_g ));
    ICE_GB masterreset_ibuf_RNIKP26_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2429),
            .GLOBALBUFFEROUTPUT(masterreset_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam masterreset_ibuf_RNIKP26_LC_12_16_3.C_ON=1'b0;
    defparam masterreset_ibuf_RNIKP26_LC_12_16_3.SEQ_MODE=4'b0000;
    defparam masterreset_ibuf_RNIKP26_LC_12_16_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 masterreset_ibuf_RNIKP26_LC_12_16_3 (
            .in0(N__3595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(masterreset_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.un3_counter_cry_1_c_LC_15_15_0 .C_ON=1'b1;
    defparam \debouncedn.un3_counter_cry_1_c_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \debouncedn.un3_counter_cry_1_c_LC_15_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debouncedn.un3_counter_cry_1_c_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__2493),
            .in2(N__2687),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\debouncedn.un3_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.un3_counter_cry_1_THRU_LUT4_0_LC_15_15_1 .C_ON=1'b1;
    defparam \debouncedn.un3_counter_cry_1_THRU_LUT4_0_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \debouncedn.un3_counter_cry_1_THRU_LUT4_0_LC_15_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debouncedn.un3_counter_cry_1_THRU_LUT4_0_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__2601),
            .in2(_gnd_net_),
            .in3(N__2519),
            .lcout(\debouncedn.un3_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\debouncedn.un3_counter_cry_1 ),
            .carryout(\debouncedn.un3_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.un3_counter_cry_2_THRU_LUT4_0_LC_15_15_2 .C_ON=1'b1;
    defparam \debouncedn.un3_counter_cry_2_THRU_LUT4_0_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \debouncedn.un3_counter_cry_2_THRU_LUT4_0_LC_15_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debouncedn.un3_counter_cry_2_THRU_LUT4_0_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__2654),
            .in2(_gnd_net_),
            .in3(N__2516),
            .lcout(\debouncedn.un3_counter_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\debouncedn.un3_counter_cry_2 ),
            .carryout(\debouncedn.un3_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_4_LC_15_15_3 .C_ON=1'b0;
    defparam \debouncedn.counter_4_LC_15_15_3 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_4_LC_15_15_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \debouncedn.counter_4_LC_15_15_3  (
            .in0(N__2476),
            .in1(N__4660),
            .in2(N__2627),
            .in3(N__2513),
            .lcout(\debouncedn.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4775),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2.C_ON=1'b0;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2 (
            .in0(N__4790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.out_RNO_1_LC_16_14_2 .C_ON=1'b0;
    defparam \debouncedn.out_RNO_1_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \debouncedn.out_RNO_1_LC_16_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \debouncedn.out_RNO_1_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__2651),
            .in2(_gnd_net_),
            .in3(N__2600),
            .lcout(),
            .ltout(\debouncedn.counter18_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.out_RNO_0_LC_16_14_3 .C_ON=1'b0;
    defparam \debouncedn.out_RNO_0_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \debouncedn.out_RNO_0_LC_16_14_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \debouncedn.out_RNO_0_LC_16_14_3  (
            .in0(N__2475),
            .in1(N__2684),
            .in2(N__2498),
            .in3(N__2494),
            .lcout(\debouncedn.out_cnv_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_1_LC_16_14_5 .C_ON=1'b0;
    defparam \debouncedn.counter_1_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_1_LC_16_14_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \debouncedn.counter_1_LC_16_14_5  (
            .in0(N__2495),
            .in1(N__2685),
            .in2(N__4666),
            .in3(N__2626),
            .lcout(\debouncedn.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4764),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_0_LC_16_15_0 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_0_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_0_LC_16_15_0 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \debounceconsolereset.counter_0_LC_16_15_0  (
            .in0(N__4587),
            .in1(_gnd_net_),
            .in2(N__2720),
            .in3(N__2811),
            .lcout(\debounceconsolereset.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4769),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_RNIBTPA2_4_LC_16_15_1 .C_ON=1'b0;
    defparam \debouncedn.counter_RNIBTPA2_4_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \debouncedn.counter_RNIBTPA2_4_LC_16_15_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \debouncedn.counter_RNIBTPA2_4_LC_16_15_1  (
            .in0(N__2652),
            .in1(N__2602),
            .in2(N__2477),
            .in3(N__4586),
            .lcout(\debouncedn.counter_RNIBTPA2Z0Z_4 ),
            .ltout(\debouncedn.counter_RNIBTPA2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_0_LC_16_15_2 .C_ON=1'b0;
    defparam \debouncedn.counter_0_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_0_LC_16_15_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \debouncedn.counter_0_LC_16_15_2  (
            .in0(N__4588),
            .in1(_gnd_net_),
            .in2(N__2690),
            .in3(N__2686),
            .lcout(\debouncedn.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4769),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_1_LC_16_15_3 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_1_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_1_LC_16_15_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \debounceconsolereset.counter_1_LC_16_15_3  (
            .in0(N__2810),
            .in1(N__2715),
            .in2(N__4663),
            .in3(N__2735),
            .lcout(\debounceconsolereset.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4769),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_RNO_1_LC_16_15_4 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNO_1_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNO_1_LC_16_15_4 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \debounceconsolereset.out_RNO_1_LC_16_15_4  (
            .in0(N__2780),
            .in1(_gnd_net_),
            .in2(N__2842),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\debounceconsolereset.counter18_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_RNO_0_LC_16_15_5 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNO_0_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNO_0_LC_16_15_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \debounceconsolereset.out_RNO_0_LC_16_15_5  (
            .in0(N__2870),
            .in1(N__2714),
            .in2(N__2663),
            .in3(N__2734),
            .lcout(\debounceconsolereset.out_cnv_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_3_LC_16_15_6 .C_ON=1'b0;
    defparam \debouncedn.counter_3_LC_16_15_6 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_3_LC_16_15_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \debouncedn.counter_3_LC_16_15_6  (
            .in0(N__2621),
            .in1(N__2660),
            .in2(N__4638),
            .in3(N__2653),
            .lcout(\debouncedn.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4769),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_2_LC_16_15_7 .C_ON=1'b0;
    defparam \debouncedn.counter_2_LC_16_15_7 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_2_LC_16_15_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \debouncedn.counter_2_LC_16_15_7  (
            .in0(N__2633),
            .in1(N__2603),
            .in2(N__4662),
            .in3(N__2622),
            .lcout(\debouncedn.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4769),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_LC_16_16_2 .C_ON=1'b0;
    defparam \debounceconsolereset.out_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.out_LC_16_16_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \debounceconsolereset.out_LC_16_16_2  (
            .in0(N__2582),
            .in1(N__2561),
            .in2(N__6107),
            .in3(N__4637),
            .lcout(debouncedconsolereset),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4776),
            .ce(),
            .sr(_gnd_net_));
    defparam lcolreg_2_LC_16_17_1.C_ON=1'b0;
    defparam lcolreg_2_LC_16_17_1.SEQ_MODE=4'b1000;
    defparam lcolreg_2_LC_16_17_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 lcolreg_2_LC_16_17_1 (
            .in0(_gnd_net_),
            .in1(N__4351),
            .in2(_gnd_net_),
            .in3(N__4488),
            .lcout(lcol3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4780),
            .ce(N__4682),
            .sr(_gnd_net_));
    defparam lcolreg_3_LC_16_17_3.C_ON=1'b0;
    defparam lcolreg_3_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam lcolreg_3_LC_16_17_3.LUT_INIT=16'b0011001111111111;
    LogicCell40 lcolreg_3_LC_16_17_3 (
            .in0(_gnd_net_),
            .in1(N__4352),
            .in2(_gnd_net_),
            .in3(N__4489),
            .lcout(lcol4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4780),
            .ce(N__4682),
            .sr(_gnd_net_));
    defparam \debounceup.un3_counter_cry_1_c_LC_17_14_0 .C_ON=1'b1;
    defparam \debounceup.un3_counter_cry_1_c_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \debounceup.un3_counter_cry_1_c_LC_17_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debounceup.un3_counter_cry_1_c_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__2940),
            .in2(N__2993),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\debounceup.un3_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.un3_counter_cry_1_THRU_LUT4_0_LC_17_14_1 .C_ON=1'b1;
    defparam \debounceup.un3_counter_cry_1_THRU_LUT4_0_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \debounceup.un3_counter_cry_1_THRU_LUT4_0_LC_17_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceup.un3_counter_cry_1_THRU_LUT4_0_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__3028),
            .in2(_gnd_net_),
            .in3(N__2756),
            .lcout(\debounceup.un3_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\debounceup.un3_counter_cry_1 ),
            .carryout(\debounceup.un3_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.un3_counter_cry_2_THRU_LUT4_0_LC_17_14_2 .C_ON=1'b1;
    defparam \debounceup.un3_counter_cry_2_THRU_LUT4_0_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \debounceup.un3_counter_cry_2_THRU_LUT4_0_LC_17_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceup.un3_counter_cry_2_THRU_LUT4_0_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__3049),
            .in2(_gnd_net_),
            .in3(N__2753),
            .lcout(\debounceup.un3_counter_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\debounceup.un3_counter_cry_2 ),
            .carryout(\debounceup.un3_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_4_LC_17_14_3 .C_ON=1'b0;
    defparam \debounceup.counter_4_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_4_LC_17_14_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \debounceup.counter_4_LC_17_14_3  (
            .in0(N__3011),
            .in1(N__4629),
            .in2(N__2969),
            .in3(N__2750),
            .lcout(\debounceup.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4760),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_3_LC_17_14_4 .C_ON=1'b0;
    defparam \debounceup.counter_3_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_3_LC_17_14_4 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \debounceup.counter_3_LC_17_14_4  (
            .in0(N__2960),
            .in1(N__2747),
            .in2(N__4665),
            .in3(N__3050),
            .lcout(\debounceup.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4760),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_2_LC_17_14_7 .C_ON=1'b0;
    defparam \debounceup.counter_2_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_2_LC_17_14_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \debounceup.counter_2_LC_17_14_7  (
            .in0(N__2741),
            .in1(N__3029),
            .in2(N__4664),
            .in3(N__2961),
            .lcout(\debounceup.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4760),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_17_15_0 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_17_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_1_c_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__2733),
            .in2(N__2719),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\debounceconsolereset.un3_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_17_15_1 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_17_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__2781),
            .in2(_gnd_net_),
            .in3(N__2696),
            .lcout(\debounceconsolereset.un3_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_1 ),
            .carryout(\debounceconsolereset.un3_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_17_15_2 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_17_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2843),
            .in3(N__2693),
            .lcout(\debounceconsolereset.un3_counter_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_2 ),
            .carryout(\debounceconsolereset.un3_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_4_LC_17_15_3 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_4_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_4_LC_17_15_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \debounceconsolereset.counter_4_LC_17_15_3  (
            .in0(N__2869),
            .in1(N__4618),
            .in2(N__2816),
            .in3(N__2873),
            .lcout(\debounceconsolereset.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4763),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_0_LC_17_15_4 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_0_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_0_LC_17_15_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \arses.clock_out_RNIR6ER_0_LC_17_15_4  (
            .in0(N__3559),
            .in1(N__3811),
            .in2(_gnd_net_),
            .in3(N__3397),
            .lcout(clock_out_RNIR6ER_0),
            .ltout(clock_out_RNIR6ER_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNINST81_4_LC_17_15_5 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_RNINST81_4_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNINST81_4_LC_17_15_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \debounceconsolereset.counter_RNINST81_4_LC_17_15_5  (
            .in0(N__2868),
            .in1(N__2837),
            .in2(N__2855),
            .in3(N__2782),
            .lcout(\debounceconsolereset.counter_RNINST81Z0Z_4 ),
            .ltout(\debounceconsolereset.counter_RNINST81Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_3_LC_17_15_6 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_3_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_3_LC_17_15_6 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \debounceconsolereset.counter_3_LC_17_15_6  (
            .in0(N__4617),
            .in1(N__2852),
            .in2(N__2846),
            .in3(N__2841),
            .lcout(\debounceconsolereset.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4763),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_2_LC_17_15_7 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_2_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_2_LC_17_15_7 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \debounceconsolereset.counter_2_LC_17_15_7  (
            .in0(N__2783),
            .in1(N__2815),
            .in2(N__2792),
            .in3(N__4619),
            .lcout(\debounceconsolereset.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4763),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.un2_counter_cry_1_c_LC_17_16_0 .C_ON=1'b1;
    defparam \arses.un2_counter_cry_1_c_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \arses.un2_counter_cry_1_c_LC_17_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \arses.un2_counter_cry_1_c_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__3254),
            .in2(N__3116),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\arses.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_2_LC_17_16_1 .C_ON=1'b1;
    defparam \arses.counter_2_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_2_LC_17_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_2_LC_17_16_1  (
            .in0(N__3411),
            .in1(N__3134),
            .in2(_gnd_net_),
            .in3(N__2762),
            .lcout(\arses.counterZ0Z_2 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_1 ),
            .carryout(\arses.un2_counter_cry_2 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_3_LC_17_16_2 .C_ON=1'b1;
    defparam \arses.counter_3_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_3_LC_17_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_3_LC_17_16_2  (
            .in0(N__3405),
            .in1(N__3146),
            .in2(_gnd_net_),
            .in3(N__2759),
            .lcout(\arses.counterZ0Z_3 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_2 ),
            .carryout(\arses.un2_counter_cry_3 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_4_LC_17_16_3 .C_ON=1'b1;
    defparam \arses.counter_4_LC_17_16_3 .SEQ_MODE=4'b1001;
    defparam \arses.counter_4_LC_17_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_4_LC_17_16_3  (
            .in0(N__3412),
            .in1(N__3266),
            .in2(_gnd_net_),
            .in3(N__2903),
            .lcout(\arses.counterZ0Z_4 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_3 ),
            .carryout(\arses.un2_counter_cry_4 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_5_LC_17_16_4 .C_ON=1'b1;
    defparam \arses.counter_5_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_5_LC_17_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_5_LC_17_16_4  (
            .in0(N__3406),
            .in1(N__3278),
            .in2(_gnd_net_),
            .in3(N__2900),
            .lcout(\arses.counterZ0Z_5 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_4 ),
            .carryout(\arses.un2_counter_cry_5 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_6_LC_17_16_5 .C_ON=1'b1;
    defparam \arses.counter_6_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_6_LC_17_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_6_LC_17_16_5  (
            .in0(N__3413),
            .in1(N__3305),
            .in2(_gnd_net_),
            .in3(N__2897),
            .lcout(\arses.counterZ0Z_6 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_5 ),
            .carryout(\arses.un2_counter_cry_6 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_7_LC_17_16_6 .C_ON=1'b1;
    defparam \arses.counter_7_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \arses.counter_7_LC_17_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_7_LC_17_16_6  (
            .in0(N__3407),
            .in1(N__3317),
            .in2(_gnd_net_),
            .in3(N__2894),
            .lcout(\arses.counterZ0Z_7 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_6 ),
            .carryout(\arses.un2_counter_cry_7 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_8_LC_17_16_7 .C_ON=1'b1;
    defparam \arses.counter_8_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \arses.counter_8_LC_17_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_8_LC_17_16_7  (
            .in0(N__3414),
            .in1(N__3292),
            .in2(_gnd_net_),
            .in3(N__2891),
            .lcout(\arses.counterZ0Z_8 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_7 ),
            .carryout(\arses.un2_counter_cry_8 ),
            .clk(N__4768),
            .ce(),
            .sr(N__4834));
    defparam \arses.counter_9_LC_17_17_0 .C_ON=1'b1;
    defparam \arses.counter_9_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \arses.counter_9_LC_17_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_9_LC_17_17_0  (
            .in0(N__3410),
            .in1(N__3200),
            .in2(_gnd_net_),
            .in3(N__2888),
            .lcout(\arses.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\arses.un2_counter_cry_9 ),
            .clk(N__4774),
            .ce(),
            .sr(N__4835));
    defparam \arses.counter_10_LC_17_17_1 .C_ON=1'b1;
    defparam \arses.counter_10_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_10_LC_17_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_10_LC_17_17_1  (
            .in0(N__3415),
            .in1(N__3215),
            .in2(_gnd_net_),
            .in3(N__2885),
            .lcout(\arses.counterZ0Z_10 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_9 ),
            .carryout(\arses.un2_counter_cry_10 ),
            .clk(N__4774),
            .ce(),
            .sr(N__4835));
    defparam \arses.counter_11_LC_17_17_2 .C_ON=1'b1;
    defparam \arses.counter_11_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_11_LC_17_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_11_LC_17_17_2  (
            .in0(N__3408),
            .in1(N__3227),
            .in2(_gnd_net_),
            .in3(N__2882),
            .lcout(\arses.counterZ0Z_11 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_10 ),
            .carryout(\arses.un2_counter_cry_11 ),
            .clk(N__4774),
            .ce(),
            .sr(N__4835));
    defparam \arses.counter_12_LC_17_17_3 .C_ON=1'b1;
    defparam \arses.counter_12_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \arses.counter_12_LC_17_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_12_LC_17_17_3  (
            .in0(N__3416),
            .in1(N__3161),
            .in2(_gnd_net_),
            .in3(N__2879),
            .lcout(\arses.counterZ0Z_12 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_11 ),
            .carryout(\arses.un2_counter_cry_12 ),
            .clk(N__4774),
            .ce(),
            .sr(N__4835));
    defparam \arses.counter_13_LC_17_17_4 .C_ON=1'b1;
    defparam \arses.counter_13_LC_17_17_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_13_LC_17_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_13_LC_17_17_4  (
            .in0(N__3409),
            .in1(N__3176),
            .in2(_gnd_net_),
            .in3(N__2876),
            .lcout(\arses.counterZ0Z_13 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_12 ),
            .carryout(\arses.un2_counter_cry_13 ),
            .clk(N__4774),
            .ce(),
            .sr(N__4835));
    defparam \arses.counter_14_LC_17_17_5 .C_ON=1'b0;
    defparam \arses.counter_14_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_14_LC_17_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_14_LC_17_17_5  (
            .in0(N__3417),
            .in1(N__3188),
            .in2(_gnd_net_),
            .in3(N__3080),
            .lcout(\arses.counterZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4774),
            .ce(),
            .sr(N__4835));
    defparam \arses.counter_1_LC_17_18_0 .C_ON=1'b0;
    defparam \arses.counter_1_LC_17_18_0 .SEQ_MODE=4'b1001;
    defparam \arses.counter_1_LC_17_18_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \arses.counter_1_LC_17_18_0  (
            .in0(N__3252),
            .in1(N__3112),
            .in2(_gnd_net_),
            .in3(N__3419),
            .lcout(\arses.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4779),
            .ce(),
            .sr(N__4836));
    defparam \dig1.leds_1_i_3_LC_18_13_0 .C_ON=1'b0;
    defparam \dig1.leds_1_i_3_LC_18_13_0 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_3_LC_18_13_0 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \dig1.leds_1_i_3_LC_18_13_0  (
            .in0(N__5729),
            .in1(N__3485),
            .in2(N__5092),
            .in3(N__3086),
            .lcout(leds_1_i_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4761),
            .ce(N__4680),
            .sr(_gnd_net_));
    defparam \debounceup.counter_RNI45V02_4_LC_18_14_2 .C_ON=1'b0;
    defparam \debounceup.counter_RNI45V02_4_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \debounceup.counter_RNI45V02_4_LC_18_14_2 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \debounceup.counter_RNI45V02_4_LC_18_14_2  (
            .in0(N__3048),
            .in1(N__3009),
            .in2(N__4639),
            .in3(N__3027),
            .lcout(\debounceup.counter_RNI45V02Z0Z_4 ),
            .ltout(\debounceup.counter_RNI45V02Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_0_LC_18_14_3 .C_ON=1'b0;
    defparam \debounceup.counter_0_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_0_LC_18_14_3 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \debounceup.counter_0_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__4595),
            .in2(N__3053),
            .in3(N__2988),
            .lcout(\debounceup.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4765),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.out_RNO_1_LC_18_14_4 .C_ON=1'b0;
    defparam \debounceup.out_RNO_1_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \debounceup.out_RNO_1_LC_18_14_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \debounceup.out_RNO_1_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__3047),
            .in2(_gnd_net_),
            .in3(N__3026),
            .lcout(),
            .ltout(\debounceup.counter18_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.out_RNO_0_LC_18_14_5 .C_ON=1'b0;
    defparam \debounceup.out_RNO_0_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \debounceup.out_RNO_0_LC_18_14_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \debounceup.out_RNO_0_LC_18_14_5  (
            .in0(N__3010),
            .in1(N__2984),
            .in2(N__2996),
            .in3(N__2941),
            .lcout(\debounceup.out_cnv_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_1_LC_18_14_6 .C_ON=1'b0;
    defparam \debounceup.counter_1_LC_18_14_6 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_1_LC_18_14_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \debounceup.counter_1_LC_18_14_6  (
            .in0(N__2942),
            .in1(N__4633),
            .in2(N__2992),
            .in3(N__2965),
            .lcout(\debounceup.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4765),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_2_LC_18_15_0 .C_ON=1'b0;
    defparam \dig1.leds_1_i_2_LC_18_15_0 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_2_LC_18_15_0 .LUT_INIT=16'b1011001110000011;
    LogicCell40 \dig1.leds_1_i_2_LC_18_15_0  (
            .in0(N__3425),
            .in1(N__3443),
            .in2(N__5737),
            .in3(N__3431),
            .lcout(leds_1_i_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4770),
            .ce(N__4681),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIA58_5_LC_18_16_2 .C_ON=1'b0;
    defparam \arses.counter_RNIA58_5_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIA58_5_LC_18_16_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \arses.counter_RNIA58_5_LC_18_16_2  (
            .in0(N__3316),
            .in1(N__3304),
            .in2(N__3293),
            .in3(N__3277),
            .lcout(),
            .ltout(\arses.un1_counterlto8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOKH_1_LC_18_16_3 .C_ON=1'b0;
    defparam \arses.counter_RNIOKH_1_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOKH_1_LC_18_16_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \arses.counter_RNIOKH_1_LC_18_16_3  (
            .in0(N__3265),
            .in1(N__3253),
            .in2(N__3230),
            .in3(N__3122),
            .lcout(),
            .ltout(\arses.un1_counterlt11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI04C4_9_LC_18_16_4 .C_ON=1'b0;
    defparam \arses.counter_RNI04C4_9_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI04C4_9_LC_18_16_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \arses.counter_RNI04C4_9_LC_18_16_4  (
            .in0(N__3226),
            .in1(N__3214),
            .in2(N__3203),
            .in3(N__3199),
            .lcout(),
            .ltout(\arses.un1_counterlt13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOS0A_14_LC_18_16_5 .C_ON=1'b0;
    defparam \arses.counter_RNIOS0A_14_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOS0A_14_LC_18_16_5 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \arses.counter_RNIOS0A_14_LC_18_16_5  (
            .in0(N__3187),
            .in1(N__3175),
            .in2(N__3164),
            .in3(N__3160),
            .lcout(\arses.counter8 ),
            .ltout(\arses.counter8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_LC_18_16_6 .C_ON=1'b0;
    defparam \arses.clock_out_LC_18_16_6 .SEQ_MODE=4'b1000;
    defparam \arses.clock_out_LC_18_16_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \arses.clock_out_LC_18_16_6  (
            .in0(N__3584),
            .in1(_gnd_net_),
            .in2(N__3149),
            .in3(N__3819),
            .lcout(slowclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4777),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI1L5_2_LC_18_17_5 .C_ON=1'b0;
    defparam \arses.counter_RNI1L5_2_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI1L5_2_LC_18_17_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \arses.counter_RNI1L5_2_LC_18_17_5  (
            .in0(N__3145),
            .in1(N__3133),
            .in2(_gnd_net_),
            .in3(N__3107),
            .lcout(\arses.un1_counterlto4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_0_LC_18_18_6 .C_ON=1'b0;
    defparam \arses.counter_0_LC_18_18_6 .SEQ_MODE=4'b1001;
    defparam \arses.counter_0_LC_18_18_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \arses.counter_0_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__3111),
            .in2(_gnd_net_),
            .in3(N__3418),
            .lcout(\arses.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4782),
            .ce(),
            .sr(N__4837));
    defparam \dig1.leds_cnst_3_1__m77_ns_LC_19_13_3 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m77_ns_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m77_ns_LC_19_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \dig1.leds_cnst_3_1__m77_ns_LC_19_13_3  (
            .in0(N__3677),
            .in1(N__3728),
            .in2(_gnd_net_),
            .in3(N__5088),
            .lcout(\dig1.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m71_LC_19_13_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m71_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m71_LC_19_13_4 .LUT_INIT=16'b0010010001000000;
    LogicCell40 \dig1.leds_cnst_3_1__m71_LC_19_13_4  (
            .in0(N__4201),
            .in1(N__5506),
            .in2(N__4490),
            .in3(N__4349),
            .lcout(\dig1.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.out_LC_19_13_5 .C_ON=1'b0;
    defparam \debouncedn.out_LC_19_13_5 .SEQ_MODE=4'b1000;
    defparam \debouncedn.out_LC_19_13_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \debouncedn.out_LC_19_13_5  (
            .in0(N__3479),
            .in1(N__3467),
            .in2(N__3509),
            .in3(N__4678),
            .lcout(debounceddn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4766),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m57_LC_19_15_3 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m57_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m57_LC_19_15_3 .LUT_INIT=16'b0011010111010010;
    LogicCell40 \dig1.leds_cnst_3_1__m57_LC_19_15_3  (
            .in0(N__4334),
            .in1(N__5496),
            .in2(N__4216),
            .in3(N__4454),
            .lcout(),
            .ltout(\dig1.N_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_15_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_15_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \dig1.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_15_4  (
            .in0(N__3437),
            .in1(N__5728),
            .in2(N__3446),
            .in3(N__5087),
            .lcout(\dig1.leds_17_i_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m60_LC_19_15_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m60_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m60_LC_19_15_5 .LUT_INIT=16'b0001110110100000;
    LogicCell40 \dig1.leds_cnst_3_1__m60_LC_19_15_5  (
            .in0(N__4333),
            .in1(N__5495),
            .in2(N__4215),
            .in3(N__4453),
            .lcout(\dig1.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m68_bm_LC_19_16_0 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m68_bm_LC_19_16_0 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m68_bm_LC_19_16_0 .LUT_INIT=16'b1001111010010010;
    LogicCell40 \dig1.leds_cnst_3_1__m68_bm_LC_19_16_0  (
            .in0(N__4466),
            .in1(N__4212),
            .in2(N__5512),
            .in3(N__4115),
            .lcout(\dig1.m68_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m68_am_LC_19_16_1 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m68_am_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m68_am_LC_19_16_1 .LUT_INIT=16'b1101000010001000;
    LogicCell40 \dig1.leds_cnst_3_1__m68_am_LC_19_16_1  (
            .in0(N__4322),
            .in1(N__5502),
            .in2(N__4217),
            .in3(N__4465),
            .lcout(\dig1.m68_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_LC_19_16_2 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_LC_19_16_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \arses.clock_out_RNIR6ER_LC_19_16_2  (
            .in0(N__3812),
            .in1(N__3583),
            .in2(_gnd_net_),
            .in3(N__3398),
            .lcout(clock_out_RNIR6ER),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam lcolreg_1_LC_19_17_6.C_ON=1'b0;
    defparam lcolreg_1_LC_19_17_6.SEQ_MODE=4'b1000;
    defparam lcolreg_1_LC_19_17_6.LUT_INIT=16'b1100110011111111;
    LogicCell40 lcolreg_1_LC_19_17_6 (
            .in0(_gnd_net_),
            .in1(N__4330),
            .in2(_gnd_net_),
            .in3(N__4471),
            .lcout(lcol2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4783),
            .ce(N__4690),
            .sr(_gnd_net_));
    defparam delayConstant_0_LC_20_11_6.C_ON=1'b0;
    defparam delayConstant_0_LC_20_11_6.SEQ_MODE=4'b1000;
    defparam delayConstant_0_LC_20_11_6.LUT_INIT=16'b0010001011011101;
    LogicCell40 delayConstant_0_LC_20_11_6 (
            .in0(N__3912),
            .in1(N__3874),
            .in2(_gnd_net_),
            .in3(N__5708),
            .lcout(delayConstantZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4762),
            .ce(),
            .sr(N__4839));
    defparam olddn_RNIM5BH1_LC_20_12_0.C_ON=1'b0;
    defparam olddn_RNIM5BH1_LC_20_12_0.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_LC_20_12_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_LC_20_12_0 (
            .in0(_gnd_net_),
            .in1(N__3907),
            .in2(_gnd_net_),
            .in3(N__3868),
            .lcout(olddn_RNIM5BHZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam oldup_RNI8NJV_LC_20_12_1.C_ON=1'b0;
    defparam oldup_RNI8NJV_LC_20_12_1.SEQ_MODE=4'b0000;
    defparam oldup_RNI8NJV_LC_20_12_1.LUT_INIT=16'b1111111101110111;
    LogicCell40 oldup_RNI8NJV_LC_20_12_1 (
            .in0(N__3585),
            .in1(N__3515),
            .in2(_gnd_net_),
            .in3(N__3690),
            .lcout(delayConstant16_i),
            .ltout(delayConstant16_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_0_c_RNO_LC_20_12_2.C_ON=1'b0;
    defparam un1_delayConstant_cry_0_c_RNO_LC_20_12_2.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_0_c_RNO_LC_20_12_2.LUT_INIT=16'b1111111100001111;
    LogicCell40 un1_delayConstant_cry_0_c_RNO_LC_20_12_2 (
            .in0(N__5712),
            .in1(_gnd_net_),
            .in2(N__3518),
            .in3(N__3867),
            .lcout(un1_delayConstant_cry_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_3_LC_20_12_3.C_ON=1'b0;
    defparam olddn_RNIM5BH1_3_LC_20_12_3.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_3_LC_20_12_3.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNIM5BH1_3_LC_20_12_3 (
            .in0(N__3869),
            .in1(_gnd_net_),
            .in2(N__3914),
            .in3(_gnd_net_),
            .lcout(olddn_RNIM5BH1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIEENH_LC_20_12_4.C_ON=1'b0;
    defparam olddn_RNIEENH_LC_20_12_4.SEQ_MODE=4'b0000;
    defparam olddn_RNIEENH_LC_20_12_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 olddn_RNIEENH_LC_20_12_4 (
            .in0(_gnd_net_),
            .in1(N__3491),
            .in2(_gnd_net_),
            .in3(N__3504),
            .lcout(olddn_RNIEENHZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam oldup_LC_20_12_5.C_ON=1'b0;
    defparam oldup_LC_20_12_5.SEQ_MODE=4'b1000;
    defparam oldup_LC_20_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 oldup_LC_20_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3691),
            .lcout(oldupZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4767),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_0_LC_20_12_6.C_ON=1'b0;
    defparam olddn_RNIM5BH1_0_LC_20_12_6.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_0_LC_20_12_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_0_LC_20_12_6 (
            .in0(_gnd_net_),
            .in1(N__3911),
            .in2(_gnd_net_),
            .in3(N__3870),
            .lcout(olddn_RNIM5BH1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_LC_20_12_7.C_ON=1'b0;
    defparam olddn_LC_20_12_7.SEQ_MODE=4'b1000;
    defparam olddn_LC_20_12_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 olddn_LC_20_12_7 (
            .in0(N__3505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(olddnZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4767),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m77_am_LC_20_13_2 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m77_am_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m77_am_LC_20_13_2 .LUT_INIT=16'b1101001110101011;
    LogicCell40 \dig1.leds_cnst_3_1__m77_am_LC_20_13_2  (
            .in0(N__4332),
            .in1(N__4172),
            .in2(N__5493),
            .in3(N__4473),
            .lcout(\dig1.m77_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.out_LC_20_13_4 .C_ON=1'b0;
    defparam \debounceup.out_LC_20_13_4 .SEQ_MODE=4'b1000;
    defparam \debounceup.out_LC_20_13_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \debounceup.out_LC_20_13_4  (
            .in0(N__3722),
            .in1(N__3692),
            .in2(N__3710),
            .in3(N__4679),
            .lcout(debouncedup),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4771),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m77_bm_LC_20_13_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m77_bm_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m77_bm_LC_20_13_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \dig1.leds_cnst_3_1__m77_bm_LC_20_13_5  (
            .in0(N__4472),
            .in1(N__4331),
            .in2(N__4197),
            .in3(N__5466),
            .lcout(\dig1.m77_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m35_LC_20_14_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m35_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m35_LC_20_14_4 .LUT_INIT=16'b0010010000001000;
    LogicCell40 \dig1.leds_cnst_3_1__m35_LC_20_14_4  (
            .in0(N__4335),
            .in1(N__5385),
            .in2(N__4050),
            .in3(N__4474),
            .lcout(\dig1.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_1_LC_20_15_3 .C_ON=1'b0;
    defparam \dig2.leds_1_i_1_LC_20_15_3 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_1_LC_20_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \dig2.leds_1_i_1_LC_20_15_3  (
            .in0(N__3830),
            .in1(N__4058),
            .in2(_gnd_net_),
            .in3(N__5779),
            .lcout(leds_1_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4781),
            .ce(N__4694),
            .sr(_gnd_net_));
    defparam lcolreg_0_LC_20_15_6.C_ON=1'b0;
    defparam lcolreg_0_LC_20_15_6.SEQ_MODE=4'b1000;
    defparam lcolreg_0_LC_20_15_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 lcolreg_0_LC_20_15_6 (
            .in0(_gnd_net_),
            .in1(N__4329),
            .in2(_gnd_net_),
            .in3(N__4470),
            .lcout(lcol1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4781),
            .ce(N__4694),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_3_LC_20_15_7 .C_ON=1'b0;
    defparam \dig2.leds_1_i_3_LC_20_15_7 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_3_LC_20_15_7 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \dig2.leds_1_i_3_LC_20_15_7  (
            .in0(N__4067),
            .in1(N__5780),
            .in2(N__5158),
            .in3(N__3632),
            .lcout(leds_1_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4781),
            .ce(N__4694),
            .sr(_gnd_net_));
    defparam col_1_LC_20_16_0.C_ON=1'b0;
    defparam col_1_LC_20_16_0.SEQ_MODE=4'b1000;
    defparam col_1_LC_20_16_0.LUT_INIT=16'b1010101011001010;
    LogicCell40 col_1_LC_20_16_0 (
            .in0(N__4311),
            .in1(N__4114),
            .in2(N__3824),
            .in3(N__3788),
            .lcout(colZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4784),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m14_LC_20_16_3 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m14_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m14_LC_20_16_3 .LUT_INIT=16'b0100011100010101;
    LogicCell40 \dig1.leds_cnst_3_1__m14_LC_20_16_3  (
            .in0(N__4047),
            .in1(N__4310),
            .in2(N__5417),
            .in3(N__4449),
            .lcout(),
            .ltout(\dig1.N_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m17_ns_LC_20_16_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m17_ns_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m17_ns_LC_20_16_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \dig1.leds_cnst_3_1__m17_ns_LC_20_16_4  (
            .in0(_gnd_net_),
            .in1(N__3779),
            .in2(N__3833),
            .in3(N__5154),
            .lcout(\dig1.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam col_0_LC_20_16_6.C_ON=1'b0;
    defparam col_0_LC_20_16_6.SEQ_MODE=4'b1000;
    defparam col_0_LC_20_16_6.LUT_INIT=16'b1010101001100110;
    LogicCell40 col_0_LC_20_16_6 (
            .in0(N__4450),
            .in1(N__3820),
            .in2(_gnd_net_),
            .in3(N__3787),
            .lcout(colZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4784),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m16_LC_20_16_7 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m16_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m16_LC_20_16_7 .LUT_INIT=16'b1010100000010010;
    LogicCell40 \dig1.leds_cnst_3_1__m16_LC_20_16_7  (
            .in0(N__4046),
            .in1(N__4309),
            .in2(N__5416),
            .in3(N__4448),
            .lcout(\dig1.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m32_am_LC_20_17_2 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m32_am_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m32_am_LC_20_17_2 .LUT_INIT=16'b1011100000001000;
    LogicCell40 \dig1.leds_cnst_3_1__m32_am_LC_20_17_2  (
            .in0(N__4052),
            .in1(N__4464),
            .in2(N__4350),
            .in3(N__5405),
            .lcout(\dig1.m32_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m32_bm_LC_20_17_7 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m32_bm_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m32_bm_LC_20_17_7 .LUT_INIT=16'b1001111010010010;
    LogicCell40 \dig1.leds_cnst_3_1__m32_bm_LC_20_17_7  (
            .in0(N__4463),
            .in1(N__4051),
            .in2(N__5418),
            .in3(N__4113),
            .lcout(\dig1.m32_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_2_LC_20_18_1 .C_ON=1'b0;
    defparam \dig2.leds_1_i_2_LC_20_18_1 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_2_LC_20_18_1 .LUT_INIT=16'b1110010001010101;
    LogicCell40 \dig2.leds_1_i_2_LC_20_18_1  (
            .in0(N__4871),
            .in1(N__3773),
            .in2(N__3767),
            .in3(N__5785),
            .lcout(leds_1_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4786),
            .ce(N__4689),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_1_LC_21_11_1.C_ON=1'b0;
    defparam olddn_RNIM5BH1_1_LC_21_11_1.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_1_LC_21_11_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_1_LC_21_11_1 (
            .in0(_gnd_net_),
            .in1(N__3904),
            .in2(_gnd_net_),
            .in3(N__3871),
            .lcout(olddn_RNIM5BH1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_4_LC_21_11_3.C_ON=1'b0;
    defparam olddn_RNIM5BH1_4_LC_21_11_3.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_4_LC_21_11_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_4_LC_21_11_3 (
            .in0(_gnd_net_),
            .in1(N__3906),
            .in2(_gnd_net_),
            .in3(N__3873),
            .lcout(olddn_RNIM5BH1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_2_LC_21_11_7.C_ON=1'b0;
    defparam olddn_RNIM5BH1_2_LC_21_11_7.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_2_LC_21_11_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_2_LC_21_11_7 (
            .in0(_gnd_net_),
            .in1(N__3905),
            .in2(_gnd_net_),
            .in3(N__3872),
            .lcout(olddn_RNIM5BH1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_0_c_LC_21_12_0.C_ON=1'b1;
    defparam un1_delayConstant_cry_0_c_LC_21_12_0.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_0_c_LC_21_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_delayConstant_cry_0_c_LC_21_12_0 (
            .in0(_gnd_net_),
            .in1(N__5697),
            .in2(N__3737),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_12_0_),
            .carryout(un1_delayConstant_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_1_LC_21_12_1.C_ON=1'b1;
    defparam delayConstant_1_LC_21_12_1.SEQ_MODE=4'b1000;
    defparam delayConstant_1_LC_21_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_1_LC_21_12_1 (
            .in0(_gnd_net_),
            .in1(N__3983),
            .in2(N__5494),
            .in3(N__3977),
            .lcout(delayConstantZ0Z_1),
            .ltout(),
            .carryin(un1_delayConstant_cry_0),
            .carryout(un1_delayConstant_cry_1),
            .clk(N__4772),
            .ce(),
            .sr(N__4840));
    defparam un1_delayConstant_cry_1_0_c_RNIJGN92_LC_21_12_2.C_ON=1'b1;
    defparam un1_delayConstant_cry_1_0_c_RNIJGN92_LC_21_12_2.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_1_0_c_RNIJGN92_LC_21_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_delayConstant_cry_1_0_c_RNIJGN92_LC_21_12_2 (
            .in0(_gnd_net_),
            .in1(N__3974),
            .in2(N__4214),
            .in3(N__3968),
            .lcout(un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92),
            .ltout(),
            .carryin(un1_delayConstant_cry_1),
            .carryout(un1_delayConstant_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_3_LC_21_12_3.C_ON=1'b1;
    defparam delayConstant_3_LC_21_12_3.SEQ_MODE=4'b1000;
    defparam delayConstant_3_LC_21_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_3_LC_21_12_3 (
            .in0(_gnd_net_),
            .in1(N__5058),
            .in2(N__3965),
            .in3(N__3956),
            .lcout(delayConstantZ0Z_3),
            .ltout(),
            .carryin(un1_delayConstant_cry_2),
            .carryout(un1_delayConstant_cry_3),
            .clk(N__4772),
            .ce(),
            .sr(N__4840));
    defparam delayConstant_4_LC_21_12_4.C_ON=1'b1;
    defparam delayConstant_4_LC_21_12_4.SEQ_MODE=4'b1000;
    defparam delayConstant_4_LC_21_12_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_4_LC_21_12_4 (
            .in0(_gnd_net_),
            .in1(N__5759),
            .in2(N__3953),
            .in3(N__3941),
            .lcout(delayConstantZ0Z_4),
            .ltout(),
            .carryin(un1_delayConstant_cry_3),
            .carryout(un1_delayConstant_cry_4),
            .clk(N__4772),
            .ce(),
            .sr(N__4840));
    defparam delayConstant_5_LC_21_12_5.C_ON=1'b1;
    defparam delayConstant_5_LC_21_12_5.SEQ_MODE=4'b1001;
    defparam delayConstant_5_LC_21_12_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_5_LC_21_12_5 (
            .in0(_gnd_net_),
            .in1(N__3938),
            .in2(N__5386),
            .in3(N__3932),
            .lcout(delayConstantZ0Z_5),
            .ltout(),
            .carryin(un1_delayConstant_cry_4),
            .carryout(un1_delayConstant_cry_5),
            .clk(N__4772),
            .ce(),
            .sr(N__4840));
    defparam un1_delayConstant_cry_5_0_c_RNIR4GA2_LC_21_12_6.C_ON=1'b1;
    defparam un1_delayConstant_cry_5_0_c_RNIR4GA2_LC_21_12_6.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_5_0_c_RNIR4GA2_LC_21_12_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_delayConstant_cry_5_0_c_RNIR4GA2_LC_21_12_6 (
            .in0(_gnd_net_),
            .in1(N__4036),
            .in2(N__3929),
            .in3(N__3917),
            .lcout(un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2),
            .ltout(),
            .carryin(un1_delayConstant_cry_5),
            .carryout(un1_delayConstant_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_7_LC_21_12_7.C_ON=1'b0;
    defparam delayConstant_7_LC_21_12_7.SEQ_MODE=4'b1000;
    defparam delayConstant_7_LC_21_12_7.LUT_INIT=16'b1000011101111000;
    LogicCell40 delayConstant_7_LC_21_12_7 (
            .in0(N__3913),
            .in1(N__3875),
            .in2(N__5153),
            .in3(N__3836),
            .lcout(delayConstantZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4772),
            .ce(),
            .sr(N__4840));
    defparam delayConstant_6_LC_21_13_6.C_ON=1'b0;
    defparam delayConstant_6_LC_21_13_6.SEQ_MODE=4'b1000;
    defparam delayConstant_6_LC_21_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_6_LC_21_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4864),
            .lcout(delayConstantZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4778),
            .ce(),
            .sr(N__4838));
    defparam delayConstant_2_LC_21_13_7.C_ON=1'b0;
    defparam delayConstant_2_LC_21_13_7.SEQ_MODE=4'b1000;
    defparam delayConstant_2_LC_21_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_2_LC_21_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4852),
            .lcout(delayConstantZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4778),
            .ce(),
            .sr(N__4838));
    defparam \dig1.leds_cnst_3_1__m41_bm_LC_21_15_2 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m41_bm_LC_21_15_2 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m41_bm_LC_21_15_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \dig1.leds_cnst_3_1__m41_bm_LC_21_15_2  (
            .in0(N__4039),
            .in1(N__4312),
            .in2(N__5406),
            .in3(N__4451),
            .lcout(\dig1.m41_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m41_am_LC_21_15_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m41_am_LC_21_15_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m41_am_LC_21_15_4 .LUT_INIT=16'b1011010111001101;
    LogicCell40 \dig1.leds_cnst_3_1__m41_am_LC_21_15_4  (
            .in0(N__4040),
            .in1(N__4313),
            .in2(N__5407),
            .in3(N__4452),
            .lcout(),
            .ltout(\dig1.m41_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m41_ns_LC_21_15_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m41_ns_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m41_ns_LC_21_15_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \dig1.leds_cnst_3_1__m41_ns_LC_21_15_5  (
            .in0(_gnd_net_),
            .in1(N__4076),
            .in2(N__4070),
            .in3(N__5147),
            .lcout(\dig1.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m2_LC_21_16_3 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m2_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m2_LC_21_16_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \dig1.leds_cnst_3_1__m2_LC_21_16_3  (
            .in0(N__4305),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4443),
            .lcout(col_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m10_ns_1_LC_21_16_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m10_ns_1_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m10_ns_1_LC_21_16_4 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \dig1.leds_cnst_3_1__m10_ns_1_LC_21_16_4  (
            .in0(N__4445),
            .in1(N__4048),
            .in2(N__5419),
            .in3(N__4306),
            .lcout(),
            .ltout(\dig1.m10_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m10_ns_LC_21_16_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m10_ns_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m10_ns_LC_21_16_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \dig1.leds_cnst_3_1__m10_ns_LC_21_16_5  (
            .in0(N__4049),
            .in1(N__4112),
            .in2(N__4061),
            .in3(N__5152),
            .lcout(\dig1.N_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m52_LC_21_16_6 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m52_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m52_LC_21_16_6 .LUT_INIT=16'b1010000110010000;
    LogicCell40 \dig1.leds_cnst_3_1__m52_LC_21_16_6  (
            .in0(N__4444),
            .in1(N__4304),
            .in2(N__4208),
            .in3(N__5489),
            .lcout(\dig1.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m24_LC_21_17_1 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m24_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m24_LC_21_17_1 .LUT_INIT=16'b0101001110001000;
    LogicCell40 \dig1.leds_cnst_3_1__m24_LC_21_17_1  (
            .in0(N__4037),
            .in1(N__4307),
            .in2(N__5414),
            .in3(N__4446),
            .lcout(\dig1.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m21_LC_21_17_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m21_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m21_LC_21_17_5 .LUT_INIT=16'b0001101110100110;
    LogicCell40 \dig1.leds_cnst_3_1__m21_LC_21_17_5  (
            .in0(N__4038),
            .in1(N__4308),
            .in2(N__5415),
            .in3(N__4447),
            .lcout(),
            .ltout(\dig1.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_21_17_6 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_21_17_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \dig1.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_21_17_6  (
            .in0(N__4880),
            .in1(N__5784),
            .in2(N__4874),
            .in3(N__5151),
            .lcout(\dig1.leds_17_i_0_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_fast_6_LC_22_11_4.C_ON=1'b0;
    defparam delayConstant_fast_6_LC_22_11_4.SEQ_MODE=4'b1000;
    defparam delayConstant_fast_6_LC_22_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_fast_6_LC_22_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4865),
            .lcout(delayConstant_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4773),
            .ce(),
            .sr(N__4841));
    defparam delayConstant_fast_2_LC_22_11_7.C_ON=1'b0;
    defparam delayConstant_fast_2_LC_22_11_7.SEQ_MODE=4'b1000;
    defparam delayConstant_fast_2_LC_22_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_fast_2_LC_22_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(delayConstant_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4773),
            .ce(),
            .sr(N__4841));
    defparam \dig1.leds_1_i_1_LC_22_15_6 .C_ON=1'b0;
    defparam \dig1.leds_1_i_1_LC_22_15_6 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_1_LC_22_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \dig1.leds_1_i_1_LC_22_15_6  (
            .in0(N__4496),
            .in1(N__4082),
            .in2(_gnd_net_),
            .in3(N__5733),
            .lcout(leds_1_i_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4785),
            .ce(N__4661),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m50_LC_22_16_1 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m50_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m50_LC_22_16_1 .LUT_INIT=16'b0001101100000111;
    LogicCell40 \dig1.leds_cnst_3_1__m50_LC_22_16_1  (
            .in0(N__4336),
            .in1(N__5508),
            .in2(N__4213),
            .in3(N__4476),
            .lcout(),
            .ltout(\dig1.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m53_ns_LC_22_16_2 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m53_ns_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m53_ns_LC_22_16_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \dig1.leds_cnst_3_1__m53_ns_LC_22_16_2  (
            .in0(_gnd_net_),
            .in1(N__5082),
            .in2(N__4505),
            .in3(N__4502),
            .lcout(\dig1.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m47_ns_1_LC_22_16_6 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m47_ns_1_LC_22_16_6 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m47_ns_1_LC_22_16_6 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \dig1.leds_cnst_3_1__m47_ns_1_LC_22_16_6  (
            .in0(N__4475),
            .in1(N__4195),
            .in2(N__5513),
            .in3(N__4337),
            .lcout(),
            .ltout(\dig1.m47_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m47_ns_LC_22_16_7 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m47_ns_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m47_ns_LC_22_16_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \dig1.leds_cnst_3_1__m47_ns_LC_22_16_7  (
            .in0(N__5083),
            .in1(N__4196),
            .in2(N__4118),
            .in3(N__4111),
            .lcout(\dig1.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_23_27_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_23_27_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_23_27_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_23_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_4_LC_27_7_5 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_4_LC_27_7_5 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_4_LC_27_7_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \arse.cpuresetoutreg_RNO_4_LC_27_7_5  (
            .in0(N__5279),
            .in1(N__5660),
            .in2(N__5639),
            .in3(N__5306),
            .lcout(\arse.g0_i_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_0_LC_27_8_0 .C_ON=1'b1;
    defparam \arse.cpuresetcount_0_LC_27_8_0 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_0_LC_27_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_0_LC_27_8_0  (
            .in0(_gnd_net_),
            .in1(N__5662),
            .in2(N__6194),
            .in3(N__6190),
            .lcout(\arse.cpuresetcountZ0Z_0 ),
            .ltout(),
            .carryin(bfn_27_8_0_),
            .carryout(\arse.un1_cpuresetcount_1_cry_0 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_1_LC_27_8_1 .C_ON=1'b1;
    defparam \arse.cpuresetcount_1_LC_27_8_1 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_1_LC_27_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_1_LC_27_8_1  (
            .in0(_gnd_net_),
            .in1(N__5282),
            .in2(_gnd_net_),
            .in3(N__4898),
            .lcout(\arse.cpuresetcountZ0Z_1 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_0 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_1 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_2_LC_27_8_2 .C_ON=1'b1;
    defparam \arse.cpuresetcount_2_LC_27_8_2 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_2_LC_27_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_2_LC_27_8_2  (
            .in0(_gnd_net_),
            .in1(N__5181),
            .in2(_gnd_net_),
            .in3(N__4895),
            .lcout(\arse.cpuresetcountZ0Z_2 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_1 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_2 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_3_LC_27_8_3 .C_ON=1'b1;
    defparam \arse.cpuresetcount_3_LC_27_8_3 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_3_LC_27_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_3_LC_27_8_3  (
            .in0(_gnd_net_),
            .in1(N__4997),
            .in2(_gnd_net_),
            .in3(N__4892),
            .lcout(\arse.cpuresetcountZ0Z_3 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_2 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_3 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_4_LC_27_8_4 .C_ON=1'b1;
    defparam \arse.cpuresetcount_4_LC_27_8_4 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_4_LC_27_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_4_LC_27_8_4  (
            .in0(_gnd_net_),
            .in1(N__5638),
            .in2(_gnd_net_),
            .in3(N__4889),
            .lcout(\arse.cpuresetcountZ0Z_4 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_3 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_4 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_5_LC_27_8_5 .C_ON=1'b1;
    defparam \arse.cpuresetcount_5_LC_27_8_5 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_5_LC_27_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_5_LC_27_8_5  (
            .in0(_gnd_net_),
            .in1(N__5309),
            .in2(_gnd_net_),
            .in3(N__4886),
            .lcout(\arse.cpuresetcountZ0Z_5 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_4 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_5 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_6_LC_27_8_6 .C_ON=1'b1;
    defparam \arse.cpuresetcount_6_LC_27_8_6 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_6_LC_27_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_6_LC_27_8_6  (
            .in0(_gnd_net_),
            .in1(N__5210),
            .in2(_gnd_net_),
            .in3(N__4883),
            .lcout(\arse.cpuresetcountZ0Z_6 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_5 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_6 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetcount_7_LC_27_8_7 .C_ON=1'b0;
    defparam \arse.cpuresetcount_7_LC_27_8_7 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_7_LC_27_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \arse.cpuresetcount_7_LC_27_8_7  (
            .in0(_gnd_net_),
            .in1(N__5020),
            .in2(_gnd_net_),
            .in3(N__5516),
            .lcout(\arse.cpuresetcountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5548));
    defparam \arse.cpuresetoutreg_RNO_2_LC_27_9_0 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_2_LC_27_9_0 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_2_LC_27_9_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \arse.cpuresetoutreg_RNO_2_LC_27_9_0  (
            .in0(N__5507),
            .in1(N__5281),
            .in2(N__5423),
            .in3(N__5307),
            .lcout(\arse.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_1_LC_28_7_0 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_1_LC_28_7_0 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_1_LC_28_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \arse.cpuresetoutreg_RNO_1_LC_28_7_0  (
            .in0(N__5016),
            .in1(N__4994),
            .in2(N__5212),
            .in3(N__5315),
            .lcout(\arse.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_RNIATKJ1_7_LC_28_7_2 .C_ON=1'b0;
    defparam \arse.cpuresetcount_RNIATKJ1_7_LC_28_7_2 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetcount_RNIATKJ1_7_LC_28_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \arse.cpuresetcount_RNIATKJ1_7_LC_28_7_2  (
            .in0(N__5015),
            .in1(N__5308),
            .in2(N__5211),
            .in3(N__5636),
            .lcout(\arse.doingseven3_6 ),
            .ltout(\arse.doingseven3_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.doingseven_RNO_0_LC_28_7_3 .C_ON=1'b0;
    defparam \arse.doingseven_RNO_0_LC_28_7_3 .SEQ_MODE=4'b0000;
    defparam \arse.doingseven_RNO_0_LC_28_7_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \arse.doingseven_RNO_0_LC_28_7_3  (
            .in0(N__4996),
            .in1(N__5258),
            .in2(N__5285),
            .in3(N__5183),
            .lcout(\arse.doingseven3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_RNIB4QP_0_LC_28_7_6 .C_ON=1'b0;
    defparam \arse.cpuresetcount_RNIB4QP_0_LC_28_7_6 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetcount_RNIB4QP_0_LC_28_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.cpuresetcount_RNIB4QP_0_LC_28_7_6  (
            .in0(_gnd_net_),
            .in1(N__5280),
            .in2(_gnd_net_),
            .in3(N__5661),
            .lcout(\arse.doingseven3_1 ),
            .ltout(\arse.doingseven3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuclkreset_RNO_0_LC_28_7_7 .C_ON=1'b0;
    defparam \arse.cpuclkreset_RNO_0_LC_28_7_7 .SEQ_MODE=4'b0000;
    defparam \arse.cpuclkreset_RNO_0_LC_28_7_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \arse.cpuclkreset_RNO_0_LC_28_7_7  (
            .in0(N__4995),
            .in1(N__5252),
            .in2(N__5246),
            .in3(N__5182),
            .lcout(\arse.doingseven4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_7_LC_28_8_0 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_7_LC_28_8_0 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_7_LC_28_8_0 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \arse.cpuresetoutreg_RNO_7_LC_28_8_0  (
            .in0(N__5243),
            .in1(N__5228),
            .in2(N__5213),
            .in3(N__5180),
            .lcout(\arse.g0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_6_LC_28_8_1 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_6_LC_28_8_1 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_6_LC_28_8_1 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \arse.cpuresetoutreg_RNO_6_LC_28_8_1  (
            .in0(N__5162),
            .in1(N__5093),
            .in2(N__5021),
            .in3(N__4993),
            .lcout(\arse.g0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_5_LC_28_8_2 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_5_LC_28_8_2 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_5_LC_28_8_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \arse.cpuresetoutreg_RNO_5_LC_28_8_2  (
            .in0(N__5786),
            .in1(N__5738),
            .in2(N__5669),
            .in3(N__5637),
            .lcout(),
            .ltout(\arse.g0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_3_LC_28_8_3 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_3_LC_28_8_3 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_3_LC_28_8_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \arse.cpuresetoutreg_RNO_3_LC_28_8_3  (
            .in0(_gnd_net_),
            .in1(N__5612),
            .in2(N__5606),
            .in3(N__5603),
            .lcout(),
            .ltout(\arse.g0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_0_LC_28_8_4 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_0_LC_28_8_4 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_0_LC_28_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \arse.cpuresetoutreg_RNO_0_LC_28_8_4  (
            .in0(N__5597),
            .in1(N__5591),
            .in2(N__5585),
            .in3(N__6189),
            .lcout(),
            .ltout(\arse.cpuresetoutreg_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_LC_28_8_5 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_LC_28_8_5 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetoutreg_LC_28_8_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \arse.cpuresetoutreg_LC_28_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5582),
            .in3(N__5575),
            .lcout(\arse.cpuresetoutregZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuresetoutregC_net ),
            .ce(),
            .sr(N__5547));
    defparam \arse.cpuclkreset_LC_29_6_6 .C_ON=1'b0;
    defparam \arse.cpuclkreset_LC_29_6_6 .SEQ_MODE=4'b1000;
    defparam \arse.cpuclkreset_LC_29_6_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \arse.cpuclkreset_LC_29_6_6  (
            .in0(N__6178),
            .in1(N__6048),
            .in2(_gnd_net_),
            .in3(N__5561),
            .lcout(\arse.cpuclkresetZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuclkresetC_net ),
            .ce(),
            .sr(N__5549));
    defparam \arse.doingseven_LC_29_7_6 .C_ON=1'b0;
    defparam \arse.doingseven_LC_29_7_6 .SEQ_MODE=4'b1000;
    defparam \arse.doingseven_LC_29_7_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \arse.doingseven_LC_29_7_6  (
            .in0(N__6179),
            .in1(N__5818),
            .in2(_gnd_net_),
            .in3(N__5555),
            .lcout(\arse.doingsevenZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.doingsevenC_net ),
            .ce(),
            .sr(N__5540));
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_4 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_4 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \debounceconsolereset.out_RNI1B6C_LC_29_8_4  (
            .in0(N__6133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debouncedconsolereset_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_0_LC_30_6_4 .C_ON=1'b0;
    defparam \arse.diveight.counter_0_LC_30_6_4 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_0_LC_30_6_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \arse.diveight.counter_0_LC_30_6_4  (
            .in0(_gnd_net_),
            .in1(N__6065),
            .in2(_gnd_net_),
            .in3(N__6039),
            .lcout(\arse.diveight.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5910),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_2_LC_30_6_5 .C_ON=1'b0;
    defparam \arse.diveight.counter_2_LC_30_6_5 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_2_LC_30_6_5 .LUT_INIT=16'b0010101010000000;
    LogicCell40 \arse.diveight.counter_2_LC_30_6_5  (
            .in0(N__6041),
            .in1(N__6010),
            .in2(N__6073),
            .in3(N__5992),
            .lcout(\arse.diveight.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5910),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_1_LC_30_6_6 .C_ON=1'b0;
    defparam \arse.diveight.counter_1_LC_30_6_6 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_1_LC_30_6_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \arse.diveight.counter_1_LC_30_6_6  (
            .in0(N__6009),
            .in1(N__6066),
            .in2(_gnd_net_),
            .in3(N__6040),
            .lcout(\arse.diveight.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5910),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.seven_LC_30_8_2 .C_ON=1'b0;
    defparam \arse.divseven.seven_LC_30_8_2 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.seven_LC_30_8_2 .LUT_INIT=16'b1110110011000100;
    LogicCell40 \arse.divseven.seven_LC_30_8_2  (
            .in0(N__5792),
            .in1(N__6232),
            .in2(N__5819),
            .in3(N__6264),
            .lcout(\arse.divseven.sevenZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5904),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_0_LC_31_6_4 .C_ON=1'b0;
    defparam \arse.diveight.dout_0_LC_31_6_4 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_0_LC_31_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.diveight.dout_0_LC_31_6_4  (
            .in0(_gnd_net_),
            .in1(N__6050),
            .in2(_gnd_net_),
            .in3(N__5991),
            .lcout(\arse.diveight.doutZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.diveight.dout_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.seven_RNO_0_LC_31_9_0 .C_ON=1'b0;
    defparam \arse.divseven.seven_RNO_0_LC_31_9_0 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.seven_RNO_0_LC_31_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.divseven.seven_RNO_0_LC_31_9_0  (
            .in0(_gnd_net_),
            .in1(N__5859),
            .in2(_gnd_net_),
            .in3(N__5952),
            .lcout(\arse.divseven.un1_counter_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_0_LC_31_9_1 .C_ON=1'b0;
    defparam \arse.divseven.counter_0_LC_31_9_1 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_0_LC_31_9_1 .LUT_INIT=16'b1000011100001111;
    LogicCell40 \arse.divseven.counter_0_LC_31_9_1  (
            .in0(N__5860),
            .in1(N__5953),
            .in2(N__6265),
            .in3(N__6230),
            .lcout(\arse.divseven.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5905),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_2_LC_31_9_2 .C_ON=1'b0;
    defparam \arse.divseven.counter_2_LC_31_9_2 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_2_LC_31_9_2 .LUT_INIT=16'b1001111111000000;
    LogicCell40 \arse.divseven.counter_2_LC_31_9_2  (
            .in0(N__6229),
            .in1(N__6257),
            .in2(N__5960),
            .in3(N__5862),
            .lcout(\arse.divseven.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5905),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_1_LC_31_9_3 .C_ON=1'b0;
    defparam \arse.divseven.counter_1_LC_31_9_3 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_1_LC_31_9_3 .LUT_INIT=16'b1011010000111100;
    LogicCell40 \arse.divseven.counter_1_LC_31_9_3  (
            .in0(N__5861),
            .in1(N__5954),
            .in2(N__6266),
            .in3(N__6231),
            .lcout(\arse.divseven.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5905),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_RNO_0_1_LC_31_9_4 .C_ON=1'b0;
    defparam \arse.divseven.dout_RNO_0_1_LC_31_9_4 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.dout_RNO_0_1_LC_31_9_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \arse.divseven.dout_RNO_0_1_LC_31_9_4  (
            .in0(N__6256),
            .in1(_gnd_net_),
            .in2(N__6233),
            .in3(_gnd_net_),
            .lcout(\arse.divseven.N_46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_RNO_0_LC_31_9_7 .C_ON=1'b0;
    defparam \arse.divseven.dout_RNO_0_LC_31_9_7 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.dout_RNO_0_LC_31_9_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \arse.divseven.dout_RNO_0_LC_31_9_7  (
            .in0(N__5858),
            .in1(N__6255),
            .in2(N__5959),
            .in3(N__6225),
            .lcout(\arse.divseven.un1_dout_2_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.apusynclatched_LC_32_4_7 .C_ON=1'b0;
    defparam \arse.apusynclatched_LC_32_4_7 .SEQ_MODE=4'b1000;
    defparam \arse.apusynclatched_LC_32_4_7 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \arse.apusynclatched_LC_32_4_7  (
            .in0(N__6153),
            .in1(N__6206),
            .in2(_gnd_net_),
            .in3(N__6132),
            .lcout(\arse.apusynclatchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.apusynclatchedC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.apuresetoutreg_LC_32_5_5 .C_ON=1'b0;
    defparam \arse.apuresetoutreg_LC_32_5_5 .SEQ_MODE=4'b1000;
    defparam \arse.apuresetoutreg_LC_32_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.apuresetoutreg_LC_32_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6140),
            .lcout(\arse.apuresetoutregZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.apuresetoutregC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_1_LC_32_6_4 .C_ON=1'b0;
    defparam \arse.diveight.dout_1_LC_32_6_4 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_1_LC_32_6_4 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \arse.diveight.dout_1_LC_32_6_4  (
            .in0(N__6074),
            .in1(N__6049),
            .in2(N__6017),
            .in3(N__5996),
            .lcout(\arse.diveight.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5912),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_1_LC_32_9_3 .C_ON=1'b0;
    defparam \arse.divseven.dout_1_LC_32_9_3 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_1_LC_32_9_3 .LUT_INIT=16'b1011110011001100;
    LogicCell40 \arse.divseven.dout_1_LC_32_9_3  (
            .in0(N__5927),
            .in1(N__5864),
            .in2(N__5969),
            .in3(N__5958),
            .lcout(\arse.divseven.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5908),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_0_LC_32_10_5 .C_ON=1'b0;
    defparam \arse.divseven.dout_0_LC_32_10_5 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_0_LC_32_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \arse.divseven.dout_0_LC_32_10_5  (
            .in0(N__5863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\arse.divseven.doutZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.divseven.dout_0C_net ),
            .ce(N__5828),
            .sr(_gnd_net_));
endmodule // top
