// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 12 2024 12:32:08

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    masterreset,
    led4,
    lcol3,
    led5,
    lcol2,
    led6,
    led2,
    lcol1,
    deldn,
    cpuclk,
    apureset,
    altreset,
    led7,
    led3,
    lcol4,
    delup,
    cpureset,
    apusync,
    PACKAGEPIN,
    led8,
    led1,
    consolereset,
    apuclk);

    input masterreset;
    output led4;
    output lcol3;
    output led5;
    output lcol2;
    output led6;
    output led2;
    output lcol1;
    input deldn;
    output cpuclk;
    output apureset;
    input altreset;
    output led7;
    output led3;
    output lcol4;
    input delup;
    output cpureset;
    input apusync;
    input PACKAGEPIN;
    output led8;
    output led1;
    input consolereset;
    output apuclk;

    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5932;
    wire N__5931;
    wire N__5930;
    wire N__5923;
    wire N__5922;
    wire N__5921;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5896;
    wire N__5895;
    wire N__5894;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5878;
    wire N__5877;
    wire N__5876;
    wire N__5869;
    wire N__5868;
    wire N__5867;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5851;
    wire N__5850;
    wire N__5849;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5833;
    wire N__5832;
    wire N__5831;
    wire N__5824;
    wire N__5823;
    wire N__5822;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5806;
    wire N__5805;
    wire N__5804;
    wire N__5797;
    wire N__5796;
    wire N__5795;
    wire N__5788;
    wire N__5787;
    wire N__5786;
    wire N__5779;
    wire N__5778;
    wire N__5777;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5761;
    wire N__5760;
    wire N__5759;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5729;
    wire N__5726;
    wire N__5725;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5704;
    wire N__5699;
    wire N__5698;
    wire N__5693;
    wire N__5690;
    wire N__5685;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5673;
    wire N__5672;
    wire N__5671;
    wire N__5668;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5656;
    wire N__5649;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5641;
    wire N__5638;
    wire N__5633;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5607;
    wire N__5606;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5589;
    wire N__5580;
    wire N__5579;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5492;
    wire N__5491;
    wire N__5490;
    wire N__5489;
    wire N__5488;
    wire N__5487;
    wire N__5484;
    wire N__5475;
    wire N__5470;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5438;
    wire N__5437;
    wire N__5436;
    wire N__5435;
    wire N__5434;
    wire N__5431;
    wire N__5422;
    wire N__5419;
    wire N__5412;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5400;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5390;
    wire N__5389;
    wire N__5388;
    wire N__5387;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5312;
    wire N__5311;
    wire N__5310;
    wire N__5309;
    wire N__5308;
    wire N__5307;
    wire N__5306;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5300;
    wire N__5299;
    wire N__5298;
    wire N__5297;
    wire N__5296;
    wire N__5295;
    wire N__5294;
    wire N__5293;
    wire N__5290;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5196;
    wire N__5195;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5187;
    wire N__5186;
    wire N__5185;
    wire N__5182;
    wire N__5173;
    wire N__5168;
    wire N__5163;
    wire N__5162;
    wire N__5161;
    wire N__5158;
    wire N__5157;
    wire N__5154;
    wire N__5153;
    wire N__5152;
    wire N__5143;
    wire N__5138;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5123;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5092;
    wire N__5089;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5075;
    wire N__5072;
    wire N__5071;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5060;
    wire N__5057;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5039;
    wire N__5032;
    wire N__5025;
    wire N__5024;
    wire N__5023;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5008;
    wire N__5001;
    wire N__4998;
    wire N__4997;
    wire N__4996;
    wire N__4995;
    wire N__4994;
    wire N__4993;
    wire N__4990;
    wire N__4983;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4979;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4961;
    wire N__4960;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4946;
    wire N__4941;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4874;
    wire N__4871;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4858;
    wire N__4851;
    wire N__4850;
    wire N__4849;
    wire N__4848;
    wire N__4845;
    wire N__4840;
    wire N__4837;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4799;
    wire N__4796;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4771;
    wire N__4764;
    wire N__4763;
    wire N__4760;
    wire N__4759;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4747;
    wire N__4740;
    wire N__4739;
    wire N__4738;
    wire N__4737;
    wire N__4736;
    wire N__4733;
    wire N__4726;
    wire N__4723;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4685;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4670;
    wire N__4669;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4650;
    wire N__4647;
    wire N__4646;
    wire N__4645;
    wire N__4644;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4596;
    wire N__4593;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4578;
    wire N__4575;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4560;
    wire N__4557;
    wire N__4556;
    wire N__4555;
    wire N__4554;
    wire N__4553;
    wire N__4552;
    wire N__4551;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4535;
    wire N__4534;
    wire N__4533;
    wire N__4524;
    wire N__4517;
    wire N__4510;
    wire N__4507;
    wire N__4502;
    wire N__4501;
    wire N__4500;
    wire N__4493;
    wire N__4486;
    wire N__4481;
    wire N__4476;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4446;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4404;
    wire N__4401;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4332;
    wire N__4329;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4317;
    wire N__4314;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4302;
    wire N__4299;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4287;
    wire N__4284;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4272;
    wire N__4269;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4254;
    wire N__4251;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4236;
    wire N__4233;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4163;
    wire N__4162;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4133;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4118;
    wire N__4113;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4064;
    wire N__4061;
    wire N__4060;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3953;
    wire N__3950;
    wire N__3949;
    wire N__3948;
    wire N__3947;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3935;
    wire N__3934;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3919;
    wire N__3918;
    wire N__3917;
    wire N__3916;
    wire N__3915;
    wire N__3914;
    wire N__3913;
    wire N__3912;
    wire N__3911;
    wire N__3910;
    wire N__3909;
    wire N__3908;
    wire N__3907;
    wire N__3906;
    wire N__3905;
    wire N__3902;
    wire N__3901;
    wire N__3900;
    wire N__3899;
    wire N__3898;
    wire N__3895;
    wire N__3890;
    wire N__3885;
    wire N__3882;
    wire N__3875;
    wire N__3872;
    wire N__3861;
    wire N__3856;
    wire N__3849;
    wire N__3844;
    wire N__3837;
    wire N__3816;
    wire N__3813;
    wire N__3812;
    wire N__3811;
    wire N__3810;
    wire N__3809;
    wire N__3806;
    wire N__3805;
    wire N__3804;
    wire N__3803;
    wire N__3798;
    wire N__3795;
    wire N__3794;
    wire N__3793;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3778;
    wire N__3773;
    wire N__3770;
    wire N__3769;
    wire N__3768;
    wire N__3767;
    wire N__3766;
    wire N__3765;
    wire N__3764;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3756;
    wire N__3755;
    wire N__3754;
    wire N__3753;
    wire N__3752;
    wire N__3751;
    wire N__3750;
    wire N__3749;
    wire N__3748;
    wire N__3747;
    wire N__3744;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3722;
    wire N__3719;
    wire N__3714;
    wire N__3709;
    wire N__3704;
    wire N__3697;
    wire N__3692;
    wire N__3685;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3629;
    wire N__3628;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3614;
    wire N__3613;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3586;
    wire N__3585;
    wire N__3584;
    wire N__3583;
    wire N__3582;
    wire N__3581;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3564;
    wire N__3559;
    wire N__3556;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3488;
    wire N__3487;
    wire N__3486;
    wire N__3485;
    wire N__3484;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3470;
    wire N__3469;
    wire N__3468;
    wire N__3467;
    wire N__3466;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3458;
    wire N__3449;
    wire N__3444;
    wire N__3441;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3403;
    wire N__3398;
    wire N__3381;
    wire N__3380;
    wire N__3379;
    wire N__3378;
    wire N__3375;
    wire N__3374;
    wire N__3373;
    wire N__3372;
    wire N__3371;
    wire N__3364;
    wire N__3361;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3343;
    wire N__3340;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3306;
    wire N__3303;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3291;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3279;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3267;
    wire N__3266;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3239;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3231;
    wire N__3228;
    wire N__3223;
    wire N__3220;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3203;
    wire N__3202;
    wire N__3201;
    wire N__3198;
    wire N__3193;
    wire N__3192;
    wire N__3189;
    wire N__3188;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3131;
    wire N__3126;
    wire N__3125;
    wire N__3124;
    wire N__3117;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3109;
    wire N__3106;
    wire N__3101;
    wire N__3096;
    wire N__3095;
    wire N__3094;
    wire N__3091;
    wire N__3086;
    wire N__3081;
    wire N__3078;
    wire N__3077;
    wire N__3076;
    wire N__3073;
    wire N__3068;
    wire N__3063;
    wire N__3062;
    wire N__3061;
    wire N__3058;
    wire N__3057;
    wire N__3054;
    wire N__3047;
    wire N__3042;
    wire N__3041;
    wire N__3040;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3028;
    wire N__3025;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3004;
    wire N__3001;
    wire N__3000;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2886;
    wire N__2885;
    wire N__2882;
    wire N__2881;
    wire N__2880;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2859;
    wire N__2856;
    wire N__2841;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2819;
    wire N__2818;
    wire N__2817;
    wire N__2816;
    wire N__2815;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2807;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2789;
    wire N__2784;
    wire N__2781;
    wire N__2780;
    wire N__2775;
    wire N__2772;
    wire N__2761;
    wire N__2758;
    wire N__2753;
    wire N__2742;
    wire N__2741;
    wire N__2740;
    wire N__2739;
    wire N__2738;
    wire N__2735;
    wire N__2734;
    wire N__2733;
    wire N__2732;
    wire N__2731;
    wire N__2730;
    wire N__2729;
    wire N__2724;
    wire N__2719;
    wire N__2716;
    wire N__2711;
    wire N__2706;
    wire N__2701;
    wire N__2696;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2658;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2646;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2622;
    wire N__2619;
    wire N__2616;
    wire N__2615;
    wire N__2614;
    wire N__2613;
    wire N__2612;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2594;
    wire N__2593;
    wire N__2590;
    wire N__2585;
    wire N__2582;
    wire N__2571;
    wire N__2562;
    wire N__2561;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2553;
    wire N__2552;
    wire N__2551;
    wire N__2550;
    wire N__2549;
    wire N__2548;
    wire N__2547;
    wire N__2544;
    wire N__2541;
    wire N__2538;
    wire N__2535;
    wire N__2522;
    wire N__2511;
    wire N__2508;
    wire N__2505;
    wire N__2502;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2454;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2424;
    wire N__2421;
    wire N__2418;
    wire N__2417;
    wire N__2412;
    wire N__2409;
    wire N__2408;
    wire N__2407;
    wire N__2404;
    wire N__2399;
    wire N__2394;
    wire N__2391;
    wire N__2388;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2376;
    wire N__2373;
    wire N__2370;
    wire N__2367;
    wire N__2364;
    wire N__2361;
    wire N__2358;
    wire N__2355;
    wire N__2352;
    wire N__2349;
    wire N__2346;
    wire N__2343;
    wire N__2340;
    wire N__2337;
    wire N__2334;
    wire N__2331;
    wire N__2328;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2316;
    wire N__2313;
    wire N__2310;
    wire N__2307;
    wire N__2304;
    wire N__2301;
    wire N__2298;
    wire N__2295;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2274;
    wire N__2271;
    wire N__2268;
    wire N__2265;
    wire N__2262;
    wire N__2259;
    wire N__2256;
    wire N__2253;
    wire N__2250;
    wire N__2247;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire \arse.un1_io_0_1_g ;
    wire \top_pll_nrtthrth.PLLOUTCORE ;
    wire \arse.divseven.io_0_D_IN_0 ;
    wire GNDG0;
    wire VCCG0;
    wire masterreset_c_i;
    wire GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO;
    wire deldn_c;
    wire leds_1_i_1;
    wire leds_1_i_3;
    wire \dig2.leds_cnst_2_cascade_ ;
    wire leds_1_i_2;
    wire olddnZ0;
    wire debounceddn;
    wire \dig2.un1_leds114_0 ;
    wire \dig2.i2_mux_cascade_ ;
    wire \dig2.leds_cnst_1 ;
    wire \dig2.m29_bm_0_cascade_ ;
    wire \dig2.m30_ns_1 ;
    wire \dig2.m23_am_0 ;
    wire \dig2.m29_am_0 ;
    wire \dig2.N_38 ;
    wire \dig2.m23_bm_0 ;
    wire \dig2.m34_am_0_cascade_ ;
    wire \dig2.m34_bm_0 ;
    wire \dig2.N_35 ;
    wire delayConstant16_i_cascade_;
    wire oldupZ0;
    wire un1_delayConstant_cry_0_c_RNOZ0;
    wire bfn_21_11_0_;
    wire olddn_RNISQ7L1Z0Z_2;
    wire un1_delayConstant_cry_0;
    wire olddn_RNISQ7L1Z0Z_0;
    wire un1_delayConstant_cry_1;
    wire olddn_RNISQ7L1Z0Z_3;
    wire un1_delayConstant_cry_2;
    wire olddn_RNISQ7L1Z0Z_1;
    wire un1_delayConstant_cry_3;
    wire olddn_RNISQ7LZ0Z1;
    wire un1_delayConstant_cry_4;
    wire olddn_RNISQ7L1Z0Z_4;
    wire un1_delayConstant_cry_5;
    wire un1_delayConstant_cry_6;
    wire delayConstant16_i;
    wire olddn_RNI1J1RZ0;
    wire delayConstantZ0Z_6;
    wire \dig2.m8_am_0_cascade_ ;
    wire \dig2.N_9 ;
    wire slowclk_0_cascade_;
    wire slowclk_0;
    wire delayConstantZ0Z_4;
    wire delayConstantZ0Z_5;
    wire \dig2.m8_bm_0 ;
    wire col_1_1;
    wire col_1_1_cascade_;
    wire \dig1.m34_am_cascade_ ;
    wire \dig1.m34_bm ;
    wire bfn_22_8_0_;
    wire \debounceconsolereset.un3_counter_cry_1 ;
    wire \debounceconsolereset.un3_counter_cry_2 ;
    wire \debounceconsolereset.un3_counter_cry_3 ;
    wire \debounceconsolereset.un3_counter_cry_2_THRU_CO ;
    wire \debounceconsolereset.un3_counter_cry_1_THRU_CO ;
    wire clock_out_RNIR6ER_0_cascade_;
    wire \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_ ;
    wire \debounceconsolereset.counter_RNINST81Z0Z_4 ;
    wire masterreset_c;
    wire slowclk;
    wire debouncedn_counter_4;
    wire debouncedn_counter_1;
    wire debouncedn_counter_0;
    wire debouncedn_counter_2;
    wire \debouncedn.out_cnvZ0Z_1 ;
    wire debouncedn_counter_3;
    wire consolereset_c;
    wire altreset_c;
    wire out_cnv_cascade_;
    wire un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2;
    wire un1_delayConstant_cry_3_0_c_RNITFZ0Z062;
    wire un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2;
    wire un1_delayConstant_cry_1_0_c_RNIP5KDZ0Z2;
    wire \dig1.m8_am_cascade_ ;
    wire \dig1.m8_bm ;
    wire \dig1.N_9_cascade_ ;
    wire \dig1.i2_mux ;
    wire \dig1.m23_bm ;
    wire \dig1.m29_bm_cascade_ ;
    wire \dig1.m23_am ;
    wire \dig1.m29_am_cascade_ ;
    wire \dig1.m30_ns_1 ;
    wire delayConstantZ0Z_0;
    wire delayConstantZ0Z_2;
    wire \dig1.leds_cnst_1 ;
    wire leds_1_i_0_1;
    wire \dig1.N_38 ;
    wire \dig1.N_35 ;
    wire leds_1_i_0_3;
    wire \dig1.un1_leds114_0 ;
    wire \dig1.leds_cnst_2 ;
    wire leds_1_i_0_2;
    wire lcol1_c;
    wire lcol2_c;
    wire lcol3_c;
    wire colZ0Z_1;
    wire colZ0Z_0;
    wire lcol4_c;
    wire clock_out_RNIR6ER_0;
    wire \INVarse.doingsevenC_net ;
    wire delayConstant_fastZ0Z_2;
    wire delayConstant_fastZ0Z_0;
    wire \arse.g0_3_cascade_ ;
    wire \arse.g0_7_cascade_ ;
    wire \arse.cpuresetoutreg_1_sqmuxa_cascade_ ;
    wire \arse.cpuresetoutregZ0 ;
    wire \INVarse.cpuresetoutregC_net ;
    wire \arses.un1_counterlto8_2_cascade_ ;
    wire \arses.un1_counterlto4_2 ;
    wire \arses.un1_counterlt11_cascade_ ;
    wire \arses.un1_counterlt13_0_cascade_ ;
    wire \arses.counterZ0Z_0 ;
    wire \arses.counterZ0Z_1 ;
    wire bfn_23_10_0_;
    wire \arses.counterZ0Z_2 ;
    wire \arses.un2_counter_cry_1 ;
    wire \arses.counterZ0Z_3 ;
    wire \arses.un2_counter_cry_2 ;
    wire \arses.counterZ0Z_4 ;
    wire \arses.un2_counter_cry_3 ;
    wire \arses.counterZ0Z_5 ;
    wire \arses.un2_counter_cry_4 ;
    wire \arses.counterZ0Z_6 ;
    wire \arses.un2_counter_cry_5 ;
    wire \arses.counterZ0Z_7 ;
    wire \arses.un2_counter_cry_6 ;
    wire \arses.counterZ0Z_8 ;
    wire \arses.un2_counter_cry_7 ;
    wire \arses.un2_counter_cry_8 ;
    wire \arses.counterZ0Z_9 ;
    wire bfn_23_11_0_;
    wire \arses.counterZ0Z_10 ;
    wire \arses.un2_counter_cry_9 ;
    wire \arses.counterZ0Z_11 ;
    wire \arses.un2_counter_cry_10 ;
    wire \arses.counterZ0Z_12 ;
    wire \arses.un2_counter_cry_11 ;
    wire \arses.counterZ0Z_13 ;
    wire \arses.un2_counter_cry_12 ;
    wire \arses.counter8 ;
    wire \arses.un2_counter_cry_13 ;
    wire \arses.counterZ0Z_14 ;
    wire masterreset_c_i_g;
    wire CONSTANT_ONE_NET;
    wire \arse.doingseven3 ;
    wire \arse.g0_i_a3_4_cascade_ ;
    wire \arse.N_6 ;
    wire \arse.doingseven3_6 ;
    wire \arse.doingseven3_1 ;
    wire \arse.doingseven3_6_cascade_ ;
    wire \arse.cpuresetcountZ0Z_0 ;
    wire bfn_24_8_0_;
    wire \arse.un1_cpuresetcount_1_cry_0 ;
    wire \arse.cpuresetcountZ0Z_2 ;
    wire \arse.un1_cpuresetcount_1_cry_1 ;
    wire \arse.un1_cpuresetcount_1_cry_2 ;
    wire \arse.un1_cpuresetcount_1_cry_3 ;
    wire \arse.un1_cpuresetcount_1_cry_4 ;
    wire \arse.un1_cpuresetcount_1_cry_5 ;
    wire \arse.un1_cpuresetcount_1_cry_6 ;
    wire \INVarse.cpuresetcount_0C_net ;
    wire delayConstantZ0Z_7;
    wire \arse.cpuresetcountZ0Z_1 ;
    wire delayConstantZ0Z_1;
    wire \arse.cpuresetcountZ0Z_7 ;
    wire \arse.g0_1 ;
    wire delayConstant_fastZ0Z_6;
    wire delayConstant_fastZ0Z_5;
    wire \arse.cpuresetcountZ0Z_6 ;
    wire \arse.cpuresetcountZ0Z_5 ;
    wire \arse.g0_4 ;
    wire delayConstant_fastZ0Z_4;
    wire delayConstantZ0Z_3;
    wire \arse.cpuresetcountZ0Z_4 ;
    wire \arse.cpuresetcountZ0Z_3 ;
    wire \arse.g0_2 ;
    wire \arse.doingsevenZ0 ;
    wire \arse.divseven.N_41_0 ;
    wire delup_c;
    wire debouncedup;
    wire PACKAGEPIN_0_c_g;
    wire out_cnv;
    wire \arse.divseven.dout_RNO_0Z0Z_0_cascade_ ;
    wire \arse.divseven.doutZ0Z_0 ;
    wire \INVarse.divseven.dout_0C_net ;
    wire \arse.divseven.counterZ0Z_1 ;
    wire \arse.divseven.sevenZ0 ;
    wire \arse.doingseven4 ;
    wire \INVarse.cpuclkresetC_net ;
    wire debouncedconsolereset_i;
    wire apusync_c;
    wire \arse.apusynclatchedZ0 ;
    wire \INVarse.apusynclatchedC_net ;
    wire \arse.diveight.counterZ0Z_0 ;
    wire \arse.diveight.counterZ0Z_1 ;
    wire \arse.diveight.doutZ0Z_1 ;
    wire \arse.cpuclkresetZ0 ;
    wire \arse.diveight.counterZ0Z_2 ;
    wire \arse.diveight.doutZ1Z_0 ;
    wire debouncedconsolereset;
    wire \arse.apuresetoutregZ0 ;
    wire \INVarse.diveight.dout_0C_net ;
    wire \arse.divseven.counterZ0Z_2 ;
    wire \arse.divseven.un1_dout_2_sqmuxa_0_o3_0 ;
    wire \arse.divseven.counterZ0Z_0 ;
    wire \arse.divseven.doutZ0Z_1 ;
    wire PLLOUTCORE_g;
    wire _gnd_net_;

    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .TEST_MODE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FILTER_RANGE=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_RELATIVE=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVR=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVQ=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVF=7'b0011111;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \top_pll_nrtthrth.top_pll_nrtthrth_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\top_pll_nrtthrth.PLLOUTCORE ),
            .REFERENCECLK(N__2337),
            .RESETB(N__3213),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF PACKAGEPIN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5959),
            .GLOBALBUFFEROUTPUT(PACKAGEPIN_0_c_g));
    IO_PAD PACKAGEPIN_ibuf_gb_io_iopad (
            .OE(N__5961),
            .DIN(N__5960),
            .DOUT(N__5959),
            .PACKAGEPIN(PACKAGEPIN));
    defparam PACKAGEPIN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam PACKAGEPIN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO PACKAGEPIN_ibuf_gb_io_preio (
            .PADOEN(N__5961),
            .PADOUT(N__5960),
            .PADIN(N__5959),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD masterreset_ibuf_iopad (
            .OE(N__5950),
            .DIN(N__5949),
            .DOUT(N__5948),
            .PACKAGEPIN(masterreset));
    defparam masterreset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam masterreset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO masterreset_ibuf_preio (
            .PADOEN(N__5950),
            .PADOUT(N__5949),
            .PADIN(N__5948),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(masterreset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led3_obuf_iopad (
            .OE(N__5941),
            .DIN(N__5940),
            .DOUT(N__5939),
            .PACKAGEPIN(led3));
    defparam led3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led3_obuf_preio (
            .PADOEN(N__5941),
            .PADOUT(N__5940),
            .PADIN(N__5939),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4044),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.divseven.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.divseven.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.divseven.io_0_iopad  (
            .OE(N__5932),
            .DIN(N__5931),
            .DOUT(N__5930),
            .PACKAGEPIN(apuclk));
    defparam \arse.divseven.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.divseven.io_0_preio  (
            .PADOEN(N__5932),
            .PADOUT(N__5931),
            .PADIN(N__5930),
            .CLOCKENABLE(),
            .DOUT1(N__5411),
            .OUTPUTENABLE(N__4415),
            .DIN0(\arse.divseven.io_0_D_IN_0 ),
            .DOUT0(N__5217),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5395));
    defparam \arse.io_1_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.io_1_iopad .PULLUP=1'b0;
    IO_PAD \arse.io_1_iopad  (
            .OE(N__5923),
            .DIN(N__5922),
            .DOUT(N__5921),
            .PACKAGEPIN(cpureset));
    defparam \arse.io_1_preio .PIN_TYPE=6'b010101;
    PRE_IO \arse.io_1_preio  (
            .PADOEN(N__5923),
            .PADOUT(N__5922),
            .PADIN(N__5921),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4206),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5400));
    IO_PAD lcol3_obuf_iopad (
            .OE(N__5914),
            .DIN(N__5913),
            .DOUT(N__5912),
            .PACKAGEPIN(lcol3));
    defparam lcol3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol3_obuf_preio (
            .PADOEN(N__5914),
            .PADOUT(N__5913),
            .PADIN(N__5912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3978),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD deldn_ibuf_iopad (
            .OE(N__5905),
            .DIN(N__5904),
            .DOUT(N__5903),
            .PACKAGEPIN(deldn));
    defparam deldn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam deldn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO deldn_ibuf_preio (
            .PADOEN(N__5905),
            .PADOUT(N__5904),
            .PADIN(N__5903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(deldn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led2_obuf_iopad (
            .OE(N__5896),
            .DIN(N__5895),
            .DOUT(N__5894),
            .PACKAGEPIN(led2));
    defparam led2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led2_obuf_preio (
            .PADOEN(N__5896),
            .PADOUT(N__5895),
            .PADIN(N__5894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3324),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delup_ibuf_iopad (
            .OE(N__5887),
            .DIN(N__5886),
            .DOUT(N__5885),
            .PACKAGEPIN(delup));
    defparam delup_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delup_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delup_ibuf_preio (
            .PADOEN(N__5887),
            .PADOUT(N__5886),
            .PADIN(N__5885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delup_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led6_obuf_iopad (
            .OE(N__5878),
            .DIN(N__5877),
            .DOUT(N__5876),
            .PACKAGEPIN(led6));
    defparam led6_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led6_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led6_obuf_preio (
            .PADOEN(N__5878),
            .PADOUT(N__5877),
            .PADIN(N__5876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led8_obuf_iopad (
            .OE(N__5869),
            .DIN(N__5868),
            .DOUT(N__5867),
            .PACKAGEPIN(led8));
    defparam led8_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led8_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led8_obuf_preio (
            .PADOEN(N__5869),
            .PADOUT(N__5868),
            .PADIN(N__5867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2283),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD altreset_ibuf_iopad (
            .OE(N__5860),
            .DIN(N__5859),
            .DOUT(N__5858),
            .PACKAGEPIN(altreset));
    defparam altreset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam altreset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO altreset_ibuf_preio (
            .PADOEN(N__5860),
            .PADOUT(N__5859),
            .PADIN(N__5858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(altreset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led4_obuf_iopad (
            .OE(N__5851),
            .DIN(N__5850),
            .DOUT(N__5849),
            .PACKAGEPIN(led4));
    defparam led4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led4_obuf_preio (
            .PADOEN(N__5851),
            .PADOUT(N__5850),
            .PADIN(N__5849),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4086),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.io_0_iopad  (
            .OE(N__5842),
            .DIN(N__5841),
            .DOUT(N__5840),
            .PACKAGEPIN(apureset));
    defparam \arse.io_0_preio .PIN_TYPE=6'b010101;
    PRE_IO \arse.io_0_preio  (
            .PADOEN(N__5842),
            .PADOUT(N__5841),
            .PADIN(N__5840),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5508),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5399));
    IO_PAD lcol4_obuf_iopad (
            .OE(N__5833),
            .DIN(N__5832),
            .DOUT(N__5831),
            .PACKAGEPIN(lcol4));
    defparam lcol4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol4_obuf_preio (
            .PADOEN(N__5833),
            .PADOUT(N__5832),
            .PADIN(N__5831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.diveight.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.diveight.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.diveight.io_0_iopad  (
            .OE(N__5824),
            .DIN(N__5823),
            .DOUT(N__5822),
            .PACKAGEPIN(cpuclk));
    defparam \arse.diveight.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.diveight.io_0_preio  (
            .PADOEN(N__5824),
            .PADOUT(N__5823),
            .PADIN(N__5822),
            .CLOCKENABLE(),
            .DOUT1(N__5628),
            .OUTPUTENABLE(N__4422),
            .DIN0(),
            .DOUT0(N__5562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5399));
    IO_PAD led5_obuf_iopad (
            .OE(N__5815),
            .DIN(N__5814),
            .DOUT(N__5813),
            .PACKAGEPIN(led5));
    defparam led5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led5_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led5_obuf_preio (
            .PADOEN(N__5815),
            .PADOUT(N__5814),
            .PADIN(N__5813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD consolereset_ibuf_iopad (
            .OE(N__5806),
            .DIN(N__5805),
            .DOUT(N__5804),
            .PACKAGEPIN(consolereset));
    defparam consolereset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam consolereset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO consolereset_ibuf_preio (
            .PADOEN(N__5806),
            .PADOUT(N__5805),
            .PADIN(N__5804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(consolereset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol2_obuf_iopad (
            .OE(N__5797),
            .DIN(N__5796),
            .DOUT(N__5795),
            .PACKAGEPIN(lcol2));
    defparam lcol2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol2_obuf_preio (
            .PADOEN(N__5797),
            .PADOUT(N__5796),
            .PADIN(N__5795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led1_obuf_iopad (
            .OE(N__5788),
            .DIN(N__5787),
            .DOUT(N__5786),
            .PACKAGEPIN(led1));
    defparam led1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led1_obuf_preio (
            .PADOEN(N__5788),
            .PADOUT(N__5787),
            .PADIN(N__5786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4393),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD apusync_ibuf_iopad (
            .OE(N__5779),
            .DIN(N__5778),
            .DOUT(N__5777),
            .PACKAGEPIN(apusync));
    defparam apusync_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam apusync_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO apusync_ibuf_preio (
            .PADOEN(N__5779),
            .PADOUT(N__5778),
            .PADIN(N__5777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(apusync_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led7_obuf_iopad (
            .OE(N__5770),
            .DIN(N__5769),
            .DOUT(N__5768),
            .PACKAGEPIN(led7));
    defparam led7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led7_obuf_preio (
            .PADOEN(N__5770),
            .PADOUT(N__5769),
            .PADIN(N__5768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2442),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol1_obuf_iopad (
            .OE(N__5761),
            .DIN(N__5760),
            .DOUT(N__5759),
            .PACKAGEPIN(lcol1));
    defparam lcol1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol1_obuf_preio (
            .PADOEN(N__5761),
            .PADOUT(N__5760),
            .PADIN(N__5759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4020),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1368 (
            .O(N__5742),
            .I(N__5739));
    LocalMux I__1367 (
            .O(N__5739),
            .I(N__5736));
    Span12Mux_v I__1366 (
            .O(N__5736),
            .I(N__5733));
    Odrv12 I__1365 (
            .O(N__5733),
            .I(apusync_c));
    InMux I__1364 (
            .O(N__5730),
            .I(N__5726));
    CascadeMux I__1363 (
            .O(N__5729),
            .I(N__5721));
    LocalMux I__1362 (
            .O(N__5726),
            .I(N__5718));
    InMux I__1361 (
            .O(N__5725),
            .I(N__5715));
    InMux I__1360 (
            .O(N__5724),
            .I(N__5712));
    InMux I__1359 (
            .O(N__5721),
            .I(N__5709));
    Span4Mux_v I__1358 (
            .O(N__5718),
            .I(N__5704));
    LocalMux I__1357 (
            .O(N__5715),
            .I(N__5704));
    LocalMux I__1356 (
            .O(N__5712),
            .I(N__5699));
    LocalMux I__1355 (
            .O(N__5709),
            .I(N__5699));
    Span4Mux_v I__1354 (
            .O(N__5704),
            .I(N__5693));
    Span4Mux_v I__1353 (
            .O(N__5699),
            .I(N__5693));
    InMux I__1352 (
            .O(N__5698),
            .I(N__5690));
    Span4Mux_h I__1351 (
            .O(N__5693),
            .I(N__5685));
    LocalMux I__1350 (
            .O(N__5690),
            .I(N__5685));
    Span4Mux_h I__1349 (
            .O(N__5685),
            .I(N__5681));
    InMux I__1348 (
            .O(N__5684),
            .I(N__5678));
    Odrv4 I__1347 (
            .O(N__5681),
            .I(\arse.apusynclatchedZ0 ));
    LocalMux I__1346 (
            .O(N__5678),
            .I(\arse.apusynclatchedZ0 ));
    CascadeMux I__1345 (
            .O(N__5673),
            .I(N__5668));
    InMux I__1344 (
            .O(N__5672),
            .I(N__5664));
    InMux I__1343 (
            .O(N__5671),
            .I(N__5661));
    InMux I__1342 (
            .O(N__5668),
            .I(N__5656));
    InMux I__1341 (
            .O(N__5667),
            .I(N__5656));
    LocalMux I__1340 (
            .O(N__5664),
            .I(\arse.diveight.counterZ0Z_0 ));
    LocalMux I__1339 (
            .O(N__5661),
            .I(\arse.diveight.counterZ0Z_0 ));
    LocalMux I__1338 (
            .O(N__5656),
            .I(\arse.diveight.counterZ0Z_0 ));
    CascadeMux I__1337 (
            .O(N__5649),
            .I(N__5645));
    CascadeMux I__1336 (
            .O(N__5648),
            .I(N__5642));
    InMux I__1335 (
            .O(N__5645),
            .I(N__5638));
    InMux I__1334 (
            .O(N__5642),
            .I(N__5633));
    InMux I__1333 (
            .O(N__5641),
            .I(N__5633));
    LocalMux I__1332 (
            .O(N__5638),
            .I(\arse.diveight.counterZ0Z_1 ));
    LocalMux I__1331 (
            .O(N__5633),
            .I(\arse.diveight.counterZ0Z_1 ));
    IoInMux I__1330 (
            .O(N__5628),
            .I(N__5625));
    LocalMux I__1329 (
            .O(N__5625),
            .I(\arse.diveight.doutZ0Z_1 ));
    InMux I__1328 (
            .O(N__5622),
            .I(N__5618));
    InMux I__1327 (
            .O(N__5621),
            .I(N__5615));
    LocalMux I__1326 (
            .O(N__5618),
            .I(N__5611));
    LocalMux I__1325 (
            .O(N__5615),
            .I(N__5608));
    InMux I__1324 (
            .O(N__5614),
            .I(N__5602));
    Span4Mux_s1_h I__1323 (
            .O(N__5611),
            .I(N__5599));
    Span4Mux_s1_h I__1322 (
            .O(N__5608),
            .I(N__5596));
    InMux I__1321 (
            .O(N__5607),
            .I(N__5589));
    InMux I__1320 (
            .O(N__5606),
            .I(N__5589));
    InMux I__1319 (
            .O(N__5605),
            .I(N__5589));
    LocalMux I__1318 (
            .O(N__5602),
            .I(\arse.cpuclkresetZ0 ));
    Odrv4 I__1317 (
            .O(N__5599),
            .I(\arse.cpuclkresetZ0 ));
    Odrv4 I__1316 (
            .O(N__5596),
            .I(\arse.cpuclkresetZ0 ));
    LocalMux I__1315 (
            .O(N__5589),
            .I(\arse.cpuclkresetZ0 ));
    InMux I__1314 (
            .O(N__5580),
            .I(N__5575));
    InMux I__1313 (
            .O(N__5579),
            .I(N__5572));
    InMux I__1312 (
            .O(N__5578),
            .I(N__5569));
    LocalMux I__1311 (
            .O(N__5575),
            .I(\arse.diveight.counterZ0Z_2 ));
    LocalMux I__1310 (
            .O(N__5572),
            .I(\arse.diveight.counterZ0Z_2 ));
    LocalMux I__1309 (
            .O(N__5569),
            .I(\arse.diveight.counterZ0Z_2 ));
    IoInMux I__1308 (
            .O(N__5562),
            .I(N__5559));
    LocalMux I__1307 (
            .O(N__5559),
            .I(\arse.diveight.doutZ1Z_0 ));
    InMux I__1306 (
            .O(N__5556),
            .I(N__5552));
    InMux I__1305 (
            .O(N__5555),
            .I(N__5549));
    LocalMux I__1304 (
            .O(N__5552),
            .I(N__5545));
    LocalMux I__1303 (
            .O(N__5549),
            .I(N__5542));
    InMux I__1302 (
            .O(N__5548),
            .I(N__5539));
    Span4Mux_v I__1301 (
            .O(N__5545),
            .I(N__5536));
    Span4Mux_s3_h I__1300 (
            .O(N__5542),
            .I(N__5531));
    LocalMux I__1299 (
            .O(N__5539),
            .I(N__5531));
    Sp12to4 I__1298 (
            .O(N__5536),
            .I(N__5528));
    Span4Mux_v I__1297 (
            .O(N__5531),
            .I(N__5525));
    Span12Mux_s10_h I__1296 (
            .O(N__5528),
            .I(N__5521));
    Sp12to4 I__1295 (
            .O(N__5525),
            .I(N__5518));
    InMux I__1294 (
            .O(N__5524),
            .I(N__5515));
    Odrv12 I__1293 (
            .O(N__5521),
            .I(debouncedconsolereset));
    Odrv12 I__1292 (
            .O(N__5518),
            .I(debouncedconsolereset));
    LocalMux I__1291 (
            .O(N__5515),
            .I(debouncedconsolereset));
    IoInMux I__1290 (
            .O(N__5508),
            .I(N__5505));
    LocalMux I__1289 (
            .O(N__5505),
            .I(\arse.apuresetoutregZ0 ));
    InMux I__1288 (
            .O(N__5502),
            .I(N__5499));
    LocalMux I__1287 (
            .O(N__5499),
            .I(N__5496));
    Span4Mux_s1_h I__1286 (
            .O(N__5496),
            .I(N__5493));
    Span4Mux_h I__1285 (
            .O(N__5493),
            .I(N__5484));
    InMux I__1284 (
            .O(N__5492),
            .I(N__5475));
    InMux I__1283 (
            .O(N__5491),
            .I(N__5475));
    InMux I__1282 (
            .O(N__5490),
            .I(N__5475));
    InMux I__1281 (
            .O(N__5489),
            .I(N__5475));
    InMux I__1280 (
            .O(N__5488),
            .I(N__5470));
    InMux I__1279 (
            .O(N__5487),
            .I(N__5470));
    Odrv4 I__1278 (
            .O(N__5484),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__1277 (
            .O(N__5475),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__1276 (
            .O(N__5470),
            .I(\arse.divseven.counterZ0Z_2 ));
    CascadeMux I__1275 (
            .O(N__5463),
            .I(N__5460));
    InMux I__1274 (
            .O(N__5460),
            .I(N__5457));
    LocalMux I__1273 (
            .O(N__5457),
            .I(N__5454));
    Span4Mux_s0_h I__1272 (
            .O(N__5454),
            .I(N__5451));
    Span4Mux_h I__1271 (
            .O(N__5451),
            .I(N__5448));
    Odrv4 I__1270 (
            .O(N__5448),
            .I(\arse.divseven.un1_dout_2_sqmuxa_0_o3_0 ));
    InMux I__1269 (
            .O(N__5445),
            .I(N__5442));
    LocalMux I__1268 (
            .O(N__5442),
            .I(N__5439));
    Span12Mux_v I__1267 (
            .O(N__5439),
            .I(N__5431));
    InMux I__1266 (
            .O(N__5438),
            .I(N__5422));
    InMux I__1265 (
            .O(N__5437),
            .I(N__5422));
    InMux I__1264 (
            .O(N__5436),
            .I(N__5422));
    InMux I__1263 (
            .O(N__5435),
            .I(N__5422));
    InMux I__1262 (
            .O(N__5434),
            .I(N__5419));
    Odrv12 I__1261 (
            .O(N__5431),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__1260 (
            .O(N__5422),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__1259 (
            .O(N__5419),
            .I(\arse.divseven.counterZ0Z_0 ));
    InMux I__1258 (
            .O(N__5412),
            .I(N__5408));
    IoInMux I__1257 (
            .O(N__5411),
            .I(N__5405));
    LocalMux I__1256 (
            .O(N__5408),
            .I(\arse.divseven.doutZ0Z_1 ));
    LocalMux I__1255 (
            .O(N__5405),
            .I(\arse.divseven.doutZ0Z_1 ));
    ClkMux I__1254 (
            .O(N__5400),
            .I(N__5358));
    ClkMux I__1253 (
            .O(N__5399),
            .I(N__5358));
    ClkMux I__1252 (
            .O(N__5398),
            .I(N__5358));
    ClkMux I__1251 (
            .O(N__5397),
            .I(N__5358));
    ClkMux I__1250 (
            .O(N__5396),
            .I(N__5358));
    ClkMux I__1249 (
            .O(N__5395),
            .I(N__5358));
    ClkMux I__1248 (
            .O(N__5394),
            .I(N__5358));
    ClkMux I__1247 (
            .O(N__5393),
            .I(N__5358));
    ClkMux I__1246 (
            .O(N__5392),
            .I(N__5358));
    ClkMux I__1245 (
            .O(N__5391),
            .I(N__5358));
    ClkMux I__1244 (
            .O(N__5390),
            .I(N__5358));
    ClkMux I__1243 (
            .O(N__5389),
            .I(N__5358));
    ClkMux I__1242 (
            .O(N__5388),
            .I(N__5358));
    ClkMux I__1241 (
            .O(N__5387),
            .I(N__5358));
    GlobalMux I__1240 (
            .O(N__5358),
            .I(N__5355));
    gio2CtrlBuf I__1239 (
            .O(N__5355),
            .I(PLLOUTCORE_g));
    CEMux I__1238 (
            .O(N__5352),
            .I(N__5349));
    LocalMux I__1237 (
            .O(N__5349),
            .I(N__5346));
    Span4Mux_h I__1236 (
            .O(N__5346),
            .I(N__5343));
    Odrv4 I__1235 (
            .O(N__5343),
            .I(\arse.divseven.N_41_0 ));
    InMux I__1234 (
            .O(N__5340),
            .I(N__5337));
    LocalMux I__1233 (
            .O(N__5337),
            .I(N__5334));
    Span12Mux_v I__1232 (
            .O(N__5334),
            .I(N__5331));
    Odrv12 I__1231 (
            .O(N__5331),
            .I(delup_c));
    InMux I__1230 (
            .O(N__5328),
            .I(N__5322));
    InMux I__1229 (
            .O(N__5327),
            .I(N__5322));
    LocalMux I__1228 (
            .O(N__5322),
            .I(N__5319));
    Odrv12 I__1227 (
            .O(N__5319),
            .I(debouncedup));
    InMux I__1226 (
            .O(N__5316),
            .I(N__5313));
    LocalMux I__1225 (
            .O(N__5313),
            .I(N__5290));
    ClkMux I__1224 (
            .O(N__5312),
            .I(N__5247));
    ClkMux I__1223 (
            .O(N__5311),
            .I(N__5247));
    ClkMux I__1222 (
            .O(N__5310),
            .I(N__5247));
    ClkMux I__1221 (
            .O(N__5309),
            .I(N__5247));
    ClkMux I__1220 (
            .O(N__5308),
            .I(N__5247));
    ClkMux I__1219 (
            .O(N__5307),
            .I(N__5247));
    ClkMux I__1218 (
            .O(N__5306),
            .I(N__5247));
    ClkMux I__1217 (
            .O(N__5305),
            .I(N__5247));
    ClkMux I__1216 (
            .O(N__5304),
            .I(N__5247));
    ClkMux I__1215 (
            .O(N__5303),
            .I(N__5247));
    ClkMux I__1214 (
            .O(N__5302),
            .I(N__5247));
    ClkMux I__1213 (
            .O(N__5301),
            .I(N__5247));
    ClkMux I__1212 (
            .O(N__5300),
            .I(N__5247));
    ClkMux I__1211 (
            .O(N__5299),
            .I(N__5247));
    ClkMux I__1210 (
            .O(N__5298),
            .I(N__5247));
    ClkMux I__1209 (
            .O(N__5297),
            .I(N__5247));
    ClkMux I__1208 (
            .O(N__5296),
            .I(N__5247));
    ClkMux I__1207 (
            .O(N__5295),
            .I(N__5247));
    ClkMux I__1206 (
            .O(N__5294),
            .I(N__5247));
    ClkMux I__1205 (
            .O(N__5293),
            .I(N__5247));
    Glb2LocalMux I__1204 (
            .O(N__5290),
            .I(N__5247));
    GlobalMux I__1203 (
            .O(N__5247),
            .I(N__5244));
    gio2CtrlBuf I__1202 (
            .O(N__5244),
            .I(PACKAGEPIN_0_c_g));
    CEMux I__1201 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__1200 (
            .O(N__5238),
            .I(N__5234));
    CEMux I__1199 (
            .O(N__5237),
            .I(N__5231));
    Span4Mux_h I__1198 (
            .O(N__5234),
            .I(N__5228));
    LocalMux I__1197 (
            .O(N__5231),
            .I(N__5225));
    Odrv4 I__1196 (
            .O(N__5228),
            .I(out_cnv));
    Odrv12 I__1195 (
            .O(N__5225),
            .I(out_cnv));
    CascadeMux I__1194 (
            .O(N__5220),
            .I(\arse.divseven.dout_RNO_0Z0Z_0_cascade_ ));
    IoInMux I__1193 (
            .O(N__5217),
            .I(N__5214));
    LocalMux I__1192 (
            .O(N__5214),
            .I(N__5211));
    IoSpan4Mux I__1191 (
            .O(N__5211),
            .I(N__5208));
    Span4Mux_s1_h I__1190 (
            .O(N__5208),
            .I(N__5204));
    InMux I__1189 (
            .O(N__5207),
            .I(N__5201));
    Odrv4 I__1188 (
            .O(N__5204),
            .I(\arse.divseven.doutZ0Z_0 ));
    LocalMux I__1187 (
            .O(N__5201),
            .I(\arse.divseven.doutZ0Z_0 ));
    CascadeMux I__1186 (
            .O(N__5196),
            .I(N__5191));
    CascadeMux I__1185 (
            .O(N__5195),
            .I(N__5188));
    CascadeMux I__1184 (
            .O(N__5194),
            .I(N__5182));
    InMux I__1183 (
            .O(N__5191),
            .I(N__5173));
    InMux I__1182 (
            .O(N__5188),
            .I(N__5173));
    InMux I__1181 (
            .O(N__5187),
            .I(N__5173));
    InMux I__1180 (
            .O(N__5186),
            .I(N__5173));
    InMux I__1179 (
            .O(N__5185),
            .I(N__5168));
    InMux I__1178 (
            .O(N__5182),
            .I(N__5168));
    LocalMux I__1177 (
            .O(N__5173),
            .I(\arse.divseven.counterZ0Z_1 ));
    LocalMux I__1176 (
            .O(N__5168),
            .I(\arse.divseven.counterZ0Z_1 ));
    CascadeMux I__1175 (
            .O(N__5163),
            .I(N__5158));
    CascadeMux I__1174 (
            .O(N__5162),
            .I(N__5154));
    InMux I__1173 (
            .O(N__5161),
            .I(N__5143));
    InMux I__1172 (
            .O(N__5158),
            .I(N__5143));
    InMux I__1171 (
            .O(N__5157),
            .I(N__5143));
    InMux I__1170 (
            .O(N__5154),
            .I(N__5143));
    InMux I__1169 (
            .O(N__5153),
            .I(N__5138));
    InMux I__1168 (
            .O(N__5152),
            .I(N__5138));
    LocalMux I__1167 (
            .O(N__5143),
            .I(\arse.divseven.sevenZ0 ));
    LocalMux I__1166 (
            .O(N__5138),
            .I(\arse.divseven.sevenZ0 ));
    InMux I__1165 (
            .O(N__5133),
            .I(N__5130));
    LocalMux I__1164 (
            .O(N__5130),
            .I(N__5127));
    Odrv12 I__1163 (
            .O(N__5127),
            .I(\arse.doingseven4 ));
    SRMux I__1162 (
            .O(N__5124),
            .I(N__5119));
    SRMux I__1161 (
            .O(N__5123),
            .I(N__5116));
    SRMux I__1160 (
            .O(N__5122),
            .I(N__5112));
    LocalMux I__1159 (
            .O(N__5119),
            .I(N__5109));
    LocalMux I__1158 (
            .O(N__5116),
            .I(N__5106));
    SRMux I__1157 (
            .O(N__5115),
            .I(N__5103));
    LocalMux I__1156 (
            .O(N__5112),
            .I(N__5100));
    Span4Mux_h I__1155 (
            .O(N__5109),
            .I(N__5097));
    Span4Mux_v I__1154 (
            .O(N__5106),
            .I(N__5092));
    LocalMux I__1153 (
            .O(N__5103),
            .I(N__5092));
    Span4Mux_v I__1152 (
            .O(N__5100),
            .I(N__5089));
    Span4Mux_v I__1151 (
            .O(N__5097),
            .I(N__5082));
    Span4Mux_h I__1150 (
            .O(N__5092),
            .I(N__5082));
    Span4Mux_v I__1149 (
            .O(N__5089),
            .I(N__5082));
    Odrv4 I__1148 (
            .O(N__5082),
            .I(debouncedconsolereset_i));
    InMux I__1147 (
            .O(N__5079),
            .I(\arse.un1_cpuresetcount_1_cry_6 ));
    CascadeMux I__1146 (
            .O(N__5076),
            .I(N__5072));
    InMux I__1145 (
            .O(N__5075),
            .I(N__5067));
    InMux I__1144 (
            .O(N__5072),
            .I(N__5064));
    InMux I__1143 (
            .O(N__5071),
            .I(N__5061));
    CascadeMux I__1142 (
            .O(N__5070),
            .I(N__5057));
    LocalMux I__1141 (
            .O(N__5067),
            .I(N__5053));
    LocalMux I__1140 (
            .O(N__5064),
            .I(N__5050));
    LocalMux I__1139 (
            .O(N__5061),
            .I(N__5047));
    InMux I__1138 (
            .O(N__5060),
            .I(N__5044));
    InMux I__1137 (
            .O(N__5057),
            .I(N__5039));
    InMux I__1136 (
            .O(N__5056),
            .I(N__5039));
    Span4Mux_h I__1135 (
            .O(N__5053),
            .I(N__5032));
    Span4Mux_h I__1134 (
            .O(N__5050),
            .I(N__5032));
    Span4Mux_h I__1133 (
            .O(N__5047),
            .I(N__5032));
    LocalMux I__1132 (
            .O(N__5044),
            .I(delayConstantZ0Z_7));
    LocalMux I__1131 (
            .O(N__5039),
            .I(delayConstantZ0Z_7));
    Odrv4 I__1130 (
            .O(N__5032),
            .I(delayConstantZ0Z_7));
    CascadeMux I__1129 (
            .O(N__5025),
            .I(N__5019));
    InMux I__1128 (
            .O(N__5024),
            .I(N__5016));
    InMux I__1127 (
            .O(N__5023),
            .I(N__5013));
    InMux I__1126 (
            .O(N__5022),
            .I(N__5008));
    InMux I__1125 (
            .O(N__5019),
            .I(N__5008));
    LocalMux I__1124 (
            .O(N__5016),
            .I(\arse.cpuresetcountZ0Z_1 ));
    LocalMux I__1123 (
            .O(N__5013),
            .I(\arse.cpuresetcountZ0Z_1 ));
    LocalMux I__1122 (
            .O(N__5008),
            .I(\arse.cpuresetcountZ0Z_1 ));
    CascadeMux I__1121 (
            .O(N__5001),
            .I(N__4998));
    InMux I__1120 (
            .O(N__4998),
            .I(N__4990));
    InMux I__1119 (
            .O(N__4997),
            .I(N__4983));
    InMux I__1118 (
            .O(N__4996),
            .I(N__4983));
    InMux I__1117 (
            .O(N__4995),
            .I(N__4983));
    InMux I__1116 (
            .O(N__4994),
            .I(N__4974));
    InMux I__1115 (
            .O(N__4993),
            .I(N__4974));
    LocalMux I__1114 (
            .O(N__4990),
            .I(N__4971));
    LocalMux I__1113 (
            .O(N__4983),
            .I(N__4968));
    InMux I__1112 (
            .O(N__4982),
            .I(N__4961));
    InMux I__1111 (
            .O(N__4981),
            .I(N__4961));
    InMux I__1110 (
            .O(N__4980),
            .I(N__4961));
    InMux I__1109 (
            .O(N__4979),
            .I(N__4956));
    LocalMux I__1108 (
            .O(N__4974),
            .I(N__4953));
    Span4Mux_h I__1107 (
            .O(N__4971),
            .I(N__4946));
    Span4Mux_v I__1106 (
            .O(N__4968),
            .I(N__4946));
    LocalMux I__1105 (
            .O(N__4961),
            .I(N__4946));
    InMux I__1104 (
            .O(N__4960),
            .I(N__4941));
    InMux I__1103 (
            .O(N__4959),
            .I(N__4941));
    LocalMux I__1102 (
            .O(N__4956),
            .I(delayConstantZ0Z_1));
    Odrv12 I__1101 (
            .O(N__4953),
            .I(delayConstantZ0Z_1));
    Odrv4 I__1100 (
            .O(N__4946),
            .I(delayConstantZ0Z_1));
    LocalMux I__1099 (
            .O(N__4941),
            .I(delayConstantZ0Z_1));
    CascadeMux I__1098 (
            .O(N__4932),
            .I(N__4926));
    InMux I__1097 (
            .O(N__4931),
            .I(N__4923));
    InMux I__1096 (
            .O(N__4930),
            .I(N__4920));
    InMux I__1095 (
            .O(N__4929),
            .I(N__4917));
    InMux I__1094 (
            .O(N__4926),
            .I(N__4914));
    LocalMux I__1093 (
            .O(N__4923),
            .I(\arse.cpuresetcountZ0Z_7 ));
    LocalMux I__1092 (
            .O(N__4920),
            .I(\arse.cpuresetcountZ0Z_7 ));
    LocalMux I__1091 (
            .O(N__4917),
            .I(\arse.cpuresetcountZ0Z_7 ));
    LocalMux I__1090 (
            .O(N__4914),
            .I(\arse.cpuresetcountZ0Z_7 ));
    InMux I__1089 (
            .O(N__4905),
            .I(N__4902));
    LocalMux I__1088 (
            .O(N__4902),
            .I(\arse.g0_1 ));
    InMux I__1087 (
            .O(N__4899),
            .I(N__4896));
    LocalMux I__1086 (
            .O(N__4896),
            .I(N__4893));
    Span4Mux_h I__1085 (
            .O(N__4893),
            .I(N__4890));
    Odrv4 I__1084 (
            .O(N__4890),
            .I(delayConstant_fastZ0Z_6));
    InMux I__1083 (
            .O(N__4887),
            .I(N__4884));
    LocalMux I__1082 (
            .O(N__4884),
            .I(N__4881));
    Span4Mux_h I__1081 (
            .O(N__4881),
            .I(N__4878));
    Odrv4 I__1080 (
            .O(N__4878),
            .I(delayConstant_fastZ0Z_5));
    CascadeMux I__1079 (
            .O(N__4875),
            .I(N__4871));
    InMux I__1078 (
            .O(N__4874),
            .I(N__4866));
    InMux I__1077 (
            .O(N__4871),
            .I(N__4863));
    InMux I__1076 (
            .O(N__4870),
            .I(N__4858));
    InMux I__1075 (
            .O(N__4869),
            .I(N__4858));
    LocalMux I__1074 (
            .O(N__4866),
            .I(\arse.cpuresetcountZ0Z_6 ));
    LocalMux I__1073 (
            .O(N__4863),
            .I(\arse.cpuresetcountZ0Z_6 ));
    LocalMux I__1072 (
            .O(N__4858),
            .I(\arse.cpuresetcountZ0Z_6 ));
    InMux I__1071 (
            .O(N__4851),
            .I(N__4845));
    InMux I__1070 (
            .O(N__4850),
            .I(N__4840));
    InMux I__1069 (
            .O(N__4849),
            .I(N__4840));
    InMux I__1068 (
            .O(N__4848),
            .I(N__4837));
    LocalMux I__1067 (
            .O(N__4845),
            .I(\arse.cpuresetcountZ0Z_5 ));
    LocalMux I__1066 (
            .O(N__4840),
            .I(\arse.cpuresetcountZ0Z_5 ));
    LocalMux I__1065 (
            .O(N__4837),
            .I(\arse.cpuresetcountZ0Z_5 ));
    InMux I__1064 (
            .O(N__4830),
            .I(N__4827));
    LocalMux I__1063 (
            .O(N__4827),
            .I(\arse.g0_4 ));
    InMux I__1062 (
            .O(N__4824),
            .I(N__4821));
    LocalMux I__1061 (
            .O(N__4821),
            .I(N__4818));
    Span4Mux_v I__1060 (
            .O(N__4818),
            .I(N__4815));
    Odrv4 I__1059 (
            .O(N__4815),
            .I(delayConstant_fastZ0Z_4));
    CascadeMux I__1058 (
            .O(N__4812),
            .I(N__4808));
    InMux I__1057 (
            .O(N__4811),
            .I(N__4805));
    InMux I__1056 (
            .O(N__4808),
            .I(N__4802));
    LocalMux I__1055 (
            .O(N__4805),
            .I(N__4796));
    LocalMux I__1054 (
            .O(N__4802),
            .I(N__4792));
    InMux I__1053 (
            .O(N__4801),
            .I(N__4789));
    InMux I__1052 (
            .O(N__4800),
            .I(N__4784));
    InMux I__1051 (
            .O(N__4799),
            .I(N__4784));
    Span4Mux_v I__1050 (
            .O(N__4796),
            .I(N__4781));
    InMux I__1049 (
            .O(N__4795),
            .I(N__4778));
    Span4Mux_v I__1048 (
            .O(N__4792),
            .I(N__4771));
    LocalMux I__1047 (
            .O(N__4789),
            .I(N__4771));
    LocalMux I__1046 (
            .O(N__4784),
            .I(N__4771));
    Odrv4 I__1045 (
            .O(N__4781),
            .I(delayConstantZ0Z_3));
    LocalMux I__1044 (
            .O(N__4778),
            .I(delayConstantZ0Z_3));
    Odrv4 I__1043 (
            .O(N__4771),
            .I(delayConstantZ0Z_3));
    CascadeMux I__1042 (
            .O(N__4764),
            .I(N__4760));
    InMux I__1041 (
            .O(N__4763),
            .I(N__4755));
    InMux I__1040 (
            .O(N__4760),
            .I(N__4752));
    InMux I__1039 (
            .O(N__4759),
            .I(N__4747));
    InMux I__1038 (
            .O(N__4758),
            .I(N__4747));
    LocalMux I__1037 (
            .O(N__4755),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1036 (
            .O(N__4752),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1035 (
            .O(N__4747),
            .I(\arse.cpuresetcountZ0Z_4 ));
    InMux I__1034 (
            .O(N__4740),
            .I(N__4733));
    InMux I__1033 (
            .O(N__4739),
            .I(N__4726));
    InMux I__1032 (
            .O(N__4738),
            .I(N__4726));
    InMux I__1031 (
            .O(N__4737),
            .I(N__4726));
    InMux I__1030 (
            .O(N__4736),
            .I(N__4723));
    LocalMux I__1029 (
            .O(N__4733),
            .I(\arse.cpuresetcountZ0Z_3 ));
    LocalMux I__1028 (
            .O(N__4726),
            .I(\arse.cpuresetcountZ0Z_3 ));
    LocalMux I__1027 (
            .O(N__4723),
            .I(\arse.cpuresetcountZ0Z_3 ));
    InMux I__1026 (
            .O(N__4716),
            .I(N__4713));
    LocalMux I__1025 (
            .O(N__4713),
            .I(\arse.g0_2 ));
    InMux I__1024 (
            .O(N__4710),
            .I(N__4706));
    InMux I__1023 (
            .O(N__4709),
            .I(N__4703));
    LocalMux I__1022 (
            .O(N__4706),
            .I(N__4700));
    LocalMux I__1021 (
            .O(N__4703),
            .I(\arse.doingsevenZ0 ));
    Odrv12 I__1020 (
            .O(N__4700),
            .I(\arse.doingsevenZ0 ));
    CascadeMux I__1019 (
            .O(N__4695),
            .I(N__4692));
    InMux I__1018 (
            .O(N__4692),
            .I(N__4689));
    LocalMux I__1017 (
            .O(N__4689),
            .I(\arse.doingseven3_6 ));
    InMux I__1016 (
            .O(N__4686),
            .I(N__4680));
    InMux I__1015 (
            .O(N__4685),
            .I(N__4680));
    LocalMux I__1014 (
            .O(N__4680),
            .I(\arse.doingseven3_1 ));
    CascadeMux I__1013 (
            .O(N__4677),
            .I(\arse.doingseven3_6_cascade_ ));
    CascadeMux I__1012 (
            .O(N__4674),
            .I(N__4671));
    InMux I__1011 (
            .O(N__4671),
            .I(N__4665));
    InMux I__1010 (
            .O(N__4670),
            .I(N__4662));
    InMux I__1009 (
            .O(N__4669),
            .I(N__4657));
    InMux I__1008 (
            .O(N__4668),
            .I(N__4657));
    LocalMux I__1007 (
            .O(N__4665),
            .I(\arse.cpuresetcountZ0Z_0 ));
    LocalMux I__1006 (
            .O(N__4662),
            .I(\arse.cpuresetcountZ0Z_0 ));
    LocalMux I__1005 (
            .O(N__4657),
            .I(\arse.cpuresetcountZ0Z_0 ));
    InMux I__1004 (
            .O(N__4650),
            .I(\arse.un1_cpuresetcount_1_cry_0 ));
    InMux I__1003 (
            .O(N__4647),
            .I(N__4639));
    InMux I__1002 (
            .O(N__4646),
            .I(N__4639));
    InMux I__1001 (
            .O(N__4645),
            .I(N__4636));
    InMux I__1000 (
            .O(N__4644),
            .I(N__4633));
    LocalMux I__999 (
            .O(N__4639),
            .I(\arse.cpuresetcountZ0Z_2 ));
    LocalMux I__998 (
            .O(N__4636),
            .I(\arse.cpuresetcountZ0Z_2 ));
    LocalMux I__997 (
            .O(N__4633),
            .I(\arse.cpuresetcountZ0Z_2 ));
    InMux I__996 (
            .O(N__4626),
            .I(\arse.un1_cpuresetcount_1_cry_1 ));
    InMux I__995 (
            .O(N__4623),
            .I(\arse.un1_cpuresetcount_1_cry_2 ));
    InMux I__994 (
            .O(N__4620),
            .I(\arse.un1_cpuresetcount_1_cry_3 ));
    InMux I__993 (
            .O(N__4617),
            .I(\arse.un1_cpuresetcount_1_cry_4 ));
    InMux I__992 (
            .O(N__4614),
            .I(\arse.un1_cpuresetcount_1_cry_5 ));
    InMux I__991 (
            .O(N__4611),
            .I(N__4607));
    InMux I__990 (
            .O(N__4610),
            .I(N__4604));
    LocalMux I__989 (
            .O(N__4607),
            .I(N__4601));
    LocalMux I__988 (
            .O(N__4604),
            .I(\arses.counterZ0Z_11 ));
    Odrv4 I__987 (
            .O(N__4601),
            .I(\arses.counterZ0Z_11 ));
    InMux I__986 (
            .O(N__4596),
            .I(\arses.un2_counter_cry_10 ));
    InMux I__985 (
            .O(N__4593),
            .I(N__4589));
    InMux I__984 (
            .O(N__4592),
            .I(N__4586));
    LocalMux I__983 (
            .O(N__4589),
            .I(N__4583));
    LocalMux I__982 (
            .O(N__4586),
            .I(\arses.counterZ0Z_12 ));
    Odrv4 I__981 (
            .O(N__4583),
            .I(\arses.counterZ0Z_12 ));
    InMux I__980 (
            .O(N__4578),
            .I(\arses.un2_counter_cry_11 ));
    InMux I__979 (
            .O(N__4575),
            .I(N__4571));
    InMux I__978 (
            .O(N__4574),
            .I(N__4568));
    LocalMux I__977 (
            .O(N__4571),
            .I(N__4565));
    LocalMux I__976 (
            .O(N__4568),
            .I(\arses.counterZ0Z_13 ));
    Odrv4 I__975 (
            .O(N__4565),
            .I(\arses.counterZ0Z_13 ));
    InMux I__974 (
            .O(N__4560),
            .I(\arses.un2_counter_cry_12 ));
    InMux I__973 (
            .O(N__4557),
            .I(N__4542));
    InMux I__972 (
            .O(N__4556),
            .I(N__4539));
    InMux I__971 (
            .O(N__4555),
            .I(N__4536));
    InMux I__970 (
            .O(N__4554),
            .I(N__4524));
    InMux I__969 (
            .O(N__4553),
            .I(N__4524));
    InMux I__968 (
            .O(N__4552),
            .I(N__4524));
    InMux I__967 (
            .O(N__4551),
            .I(N__4524));
    InMux I__966 (
            .O(N__4550),
            .I(N__4517));
    InMux I__965 (
            .O(N__4549),
            .I(N__4517));
    InMux I__964 (
            .O(N__4548),
            .I(N__4517));
    InMux I__963 (
            .O(N__4547),
            .I(N__4510));
    InMux I__962 (
            .O(N__4546),
            .I(N__4510));
    InMux I__961 (
            .O(N__4545),
            .I(N__4510));
    LocalMux I__960 (
            .O(N__4542),
            .I(N__4507));
    LocalMux I__959 (
            .O(N__4539),
            .I(N__4502));
    LocalMux I__958 (
            .O(N__4536),
            .I(N__4502));
    InMux I__957 (
            .O(N__4535),
            .I(N__4493));
    InMux I__956 (
            .O(N__4534),
            .I(N__4493));
    InMux I__955 (
            .O(N__4533),
            .I(N__4493));
    LocalMux I__954 (
            .O(N__4524),
            .I(N__4486));
    LocalMux I__953 (
            .O(N__4517),
            .I(N__4486));
    LocalMux I__952 (
            .O(N__4510),
            .I(N__4486));
    Span4Mux_h I__951 (
            .O(N__4507),
            .I(N__4481));
    Span4Mux_v I__950 (
            .O(N__4502),
            .I(N__4481));
    InMux I__949 (
            .O(N__4501),
            .I(N__4476));
    InMux I__948 (
            .O(N__4500),
            .I(N__4476));
    LocalMux I__947 (
            .O(N__4493),
            .I(\arses.counter8 ));
    Odrv4 I__946 (
            .O(N__4486),
            .I(\arses.counter8 ));
    Odrv4 I__945 (
            .O(N__4481),
            .I(\arses.counter8 ));
    LocalMux I__944 (
            .O(N__4476),
            .I(\arses.counter8 ));
    InMux I__943 (
            .O(N__4467),
            .I(\arses.un2_counter_cry_13 ));
    InMux I__942 (
            .O(N__4464),
            .I(N__4461));
    LocalMux I__941 (
            .O(N__4461),
            .I(N__4457));
    InMux I__940 (
            .O(N__4460),
            .I(N__4454));
    Span4Mux_h I__939 (
            .O(N__4457),
            .I(N__4451));
    LocalMux I__938 (
            .O(N__4454),
            .I(\arses.counterZ0Z_14 ));
    Odrv4 I__937 (
            .O(N__4451),
            .I(\arses.counterZ0Z_14 ));
    SRMux I__936 (
            .O(N__4446),
            .I(N__4428));
    SRMux I__935 (
            .O(N__4445),
            .I(N__4428));
    SRMux I__934 (
            .O(N__4444),
            .I(N__4428));
    SRMux I__933 (
            .O(N__4443),
            .I(N__4428));
    SRMux I__932 (
            .O(N__4442),
            .I(N__4428));
    SRMux I__931 (
            .O(N__4441),
            .I(N__4428));
    GlobalMux I__930 (
            .O(N__4428),
            .I(N__4425));
    gio2CtrlBuf I__929 (
            .O(N__4425),
            .I(masterreset_c_i_g));
    IoInMux I__928 (
            .O(N__4422),
            .I(N__4419));
    LocalMux I__927 (
            .O(N__4419),
            .I(N__4416));
    IoSpan4Mux I__926 (
            .O(N__4416),
            .I(N__4412));
    IoInMux I__925 (
            .O(N__4415),
            .I(N__4409));
    IoSpan4Mux I__924 (
            .O(N__4412),
            .I(N__4404));
    LocalMux I__923 (
            .O(N__4409),
            .I(N__4404));
    Span4Mux_s2_h I__922 (
            .O(N__4404),
            .I(N__4401));
    Span4Mux_h I__921 (
            .O(N__4401),
            .I(N__4397));
    IoInMux I__920 (
            .O(N__4400),
            .I(N__4394));
    Sp12to4 I__919 (
            .O(N__4397),
            .I(N__4390));
    LocalMux I__918 (
            .O(N__4394),
            .I(N__4387));
    IoInMux I__917 (
            .O(N__4393),
            .I(N__4384));
    Span12Mux_v I__916 (
            .O(N__4390),
            .I(N__4381));
    Span4Mux_s1_v I__915 (
            .O(N__4387),
            .I(N__4378));
    LocalMux I__914 (
            .O(N__4384),
            .I(N__4375));
    Span12Mux_v I__913 (
            .O(N__4381),
            .I(N__4372));
    Span4Mux_h I__912 (
            .O(N__4378),
            .I(N__4369));
    Span12Mux_s1_v I__911 (
            .O(N__4375),
            .I(N__4366));
    Odrv12 I__910 (
            .O(N__4372),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__909 (
            .O(N__4369),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__908 (
            .O(N__4366),
            .I(CONSTANT_ONE_NET));
    InMux I__907 (
            .O(N__4359),
            .I(N__4356));
    LocalMux I__906 (
            .O(N__4356),
            .I(\arse.doingseven3 ));
    CascadeMux I__905 (
            .O(N__4353),
            .I(\arse.g0_i_a3_4_cascade_ ));
    InMux I__904 (
            .O(N__4350),
            .I(N__4347));
    LocalMux I__903 (
            .O(N__4347),
            .I(\arse.N_6 ));
    InMux I__902 (
            .O(N__4344),
            .I(N__4340));
    InMux I__901 (
            .O(N__4343),
            .I(N__4337));
    LocalMux I__900 (
            .O(N__4340),
            .I(\arses.counterZ0Z_3 ));
    LocalMux I__899 (
            .O(N__4337),
            .I(\arses.counterZ0Z_3 ));
    InMux I__898 (
            .O(N__4332),
            .I(\arses.un2_counter_cry_2 ));
    InMux I__897 (
            .O(N__4329),
            .I(N__4325));
    InMux I__896 (
            .O(N__4328),
            .I(N__4322));
    LocalMux I__895 (
            .O(N__4325),
            .I(\arses.counterZ0Z_4 ));
    LocalMux I__894 (
            .O(N__4322),
            .I(\arses.counterZ0Z_4 ));
    InMux I__893 (
            .O(N__4317),
            .I(\arses.un2_counter_cry_3 ));
    InMux I__892 (
            .O(N__4314),
            .I(N__4310));
    InMux I__891 (
            .O(N__4313),
            .I(N__4307));
    LocalMux I__890 (
            .O(N__4310),
            .I(\arses.counterZ0Z_5 ));
    LocalMux I__889 (
            .O(N__4307),
            .I(\arses.counterZ0Z_5 ));
    InMux I__888 (
            .O(N__4302),
            .I(\arses.un2_counter_cry_4 ));
    InMux I__887 (
            .O(N__4299),
            .I(N__4295));
    InMux I__886 (
            .O(N__4298),
            .I(N__4292));
    LocalMux I__885 (
            .O(N__4295),
            .I(\arses.counterZ0Z_6 ));
    LocalMux I__884 (
            .O(N__4292),
            .I(\arses.counterZ0Z_6 ));
    InMux I__883 (
            .O(N__4287),
            .I(\arses.un2_counter_cry_5 ));
    InMux I__882 (
            .O(N__4284),
            .I(N__4280));
    InMux I__881 (
            .O(N__4283),
            .I(N__4277));
    LocalMux I__880 (
            .O(N__4280),
            .I(\arses.counterZ0Z_7 ));
    LocalMux I__879 (
            .O(N__4277),
            .I(\arses.counterZ0Z_7 ));
    InMux I__878 (
            .O(N__4272),
            .I(\arses.un2_counter_cry_6 ));
    CascadeMux I__877 (
            .O(N__4269),
            .I(N__4265));
    InMux I__876 (
            .O(N__4268),
            .I(N__4262));
    InMux I__875 (
            .O(N__4265),
            .I(N__4259));
    LocalMux I__874 (
            .O(N__4262),
            .I(\arses.counterZ0Z_8 ));
    LocalMux I__873 (
            .O(N__4259),
            .I(\arses.counterZ0Z_8 ));
    InMux I__872 (
            .O(N__4254),
            .I(\arses.un2_counter_cry_7 ));
    InMux I__871 (
            .O(N__4251),
            .I(N__4247));
    InMux I__870 (
            .O(N__4250),
            .I(N__4244));
    LocalMux I__869 (
            .O(N__4247),
            .I(N__4241));
    LocalMux I__868 (
            .O(N__4244),
            .I(\arses.counterZ0Z_9 ));
    Odrv4 I__867 (
            .O(N__4241),
            .I(\arses.counterZ0Z_9 ));
    InMux I__866 (
            .O(N__4236),
            .I(bfn_23_11_0_));
    InMux I__865 (
            .O(N__4233),
            .I(N__4229));
    InMux I__864 (
            .O(N__4232),
            .I(N__4226));
    LocalMux I__863 (
            .O(N__4229),
            .I(N__4223));
    LocalMux I__862 (
            .O(N__4226),
            .I(\arses.counterZ0Z_10 ));
    Odrv4 I__861 (
            .O(N__4223),
            .I(\arses.counterZ0Z_10 ));
    InMux I__860 (
            .O(N__4218),
            .I(\arses.un2_counter_cry_9 ));
    CascadeMux I__859 (
            .O(N__4215),
            .I(\arse.g0_3_cascade_ ));
    CascadeMux I__858 (
            .O(N__4212),
            .I(\arse.g0_7_cascade_ ));
    CascadeMux I__857 (
            .O(N__4209),
            .I(\arse.cpuresetoutreg_1_sqmuxa_cascade_ ));
    IoInMux I__856 (
            .O(N__4206),
            .I(N__4203));
    LocalMux I__855 (
            .O(N__4203),
            .I(N__4200));
    Span4Mux_s0_h I__854 (
            .O(N__4200),
            .I(N__4197));
    Span4Mux_h I__853 (
            .O(N__4197),
            .I(N__4193));
    InMux I__852 (
            .O(N__4196),
            .I(N__4190));
    Span4Mux_h I__851 (
            .O(N__4193),
            .I(N__4187));
    LocalMux I__850 (
            .O(N__4190),
            .I(\arse.cpuresetoutregZ0 ));
    Odrv4 I__849 (
            .O(N__4187),
            .I(\arse.cpuresetoutregZ0 ));
    CascadeMux I__848 (
            .O(N__4182),
            .I(\arses.un1_counterlto8_2_cascade_ ));
    InMux I__847 (
            .O(N__4179),
            .I(N__4176));
    LocalMux I__846 (
            .O(N__4176),
            .I(\arses.un1_counterlto4_2 ));
    CascadeMux I__845 (
            .O(N__4173),
            .I(\arses.un1_counterlt11_cascade_ ));
    CascadeMux I__844 (
            .O(N__4170),
            .I(\arses.un1_counterlt13_0_cascade_ ));
    InMux I__843 (
            .O(N__4167),
            .I(N__4164));
    LocalMux I__842 (
            .O(N__4164),
            .I(N__4158));
    InMux I__841 (
            .O(N__4163),
            .I(N__4155));
    InMux I__840 (
            .O(N__4162),
            .I(N__4152));
    InMux I__839 (
            .O(N__4161),
            .I(N__4149));
    Odrv4 I__838 (
            .O(N__4158),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__837 (
            .O(N__4155),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__836 (
            .O(N__4152),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__835 (
            .O(N__4149),
            .I(\arses.counterZ0Z_0 ));
    CascadeMux I__834 (
            .O(N__4140),
            .I(N__4137));
    InMux I__833 (
            .O(N__4137),
            .I(N__4134));
    LocalMux I__832 (
            .O(N__4134),
            .I(N__4129));
    InMux I__831 (
            .O(N__4133),
            .I(N__4126));
    InMux I__830 (
            .O(N__4132),
            .I(N__4123));
    Span4Mux_v I__829 (
            .O(N__4129),
            .I(N__4118));
    LocalMux I__828 (
            .O(N__4126),
            .I(N__4118));
    LocalMux I__827 (
            .O(N__4123),
            .I(\arses.counterZ0Z_1 ));
    Odrv4 I__826 (
            .O(N__4118),
            .I(\arses.counterZ0Z_1 ));
    InMux I__825 (
            .O(N__4113),
            .I(N__4109));
    InMux I__824 (
            .O(N__4112),
            .I(N__4106));
    LocalMux I__823 (
            .O(N__4109),
            .I(\arses.counterZ0Z_2 ));
    LocalMux I__822 (
            .O(N__4106),
            .I(\arses.counterZ0Z_2 ));
    InMux I__821 (
            .O(N__4101),
            .I(\arses.un2_counter_cry_1 ));
    InMux I__820 (
            .O(N__4098),
            .I(N__4095));
    LocalMux I__819 (
            .O(N__4095),
            .I(\dig1.N_38 ));
    InMux I__818 (
            .O(N__4092),
            .I(N__4089));
    LocalMux I__817 (
            .O(N__4089),
            .I(\dig1.N_35 ));
    IoInMux I__816 (
            .O(N__4086),
            .I(N__4083));
    LocalMux I__815 (
            .O(N__4083),
            .I(N__4080));
    IoSpan4Mux I__814 (
            .O(N__4080),
            .I(N__4077));
    Sp12to4 I__813 (
            .O(N__4077),
            .I(N__4074));
    Span12Mux_s6_v I__812 (
            .O(N__4074),
            .I(N__4071));
    Span12Mux_h I__811 (
            .O(N__4071),
            .I(N__4068));
    Odrv12 I__810 (
            .O(N__4068),
            .I(leds_1_i_0_3));
    CascadeMux I__809 (
            .O(N__4065),
            .I(N__4061));
    InMux I__808 (
            .O(N__4064),
            .I(N__4053));
    InMux I__807 (
            .O(N__4061),
            .I(N__4053));
    InMux I__806 (
            .O(N__4060),
            .I(N__4053));
    LocalMux I__805 (
            .O(N__4053),
            .I(\dig1.un1_leds114_0 ));
    InMux I__804 (
            .O(N__4050),
            .I(N__4047));
    LocalMux I__803 (
            .O(N__4047),
            .I(\dig1.leds_cnst_2 ));
    IoInMux I__802 (
            .O(N__4044),
            .I(N__4041));
    LocalMux I__801 (
            .O(N__4041),
            .I(N__4038));
    Span4Mux_s1_v I__800 (
            .O(N__4038),
            .I(N__4035));
    Span4Mux_v I__799 (
            .O(N__4035),
            .I(N__4032));
    Sp12to4 I__798 (
            .O(N__4032),
            .I(N__4029));
    Span12Mux_h I__797 (
            .O(N__4029),
            .I(N__4026));
    Span12Mux_v I__796 (
            .O(N__4026),
            .I(N__4023));
    Odrv12 I__795 (
            .O(N__4023),
            .I(leds_1_i_0_2));
    IoInMux I__794 (
            .O(N__4020),
            .I(N__4017));
    LocalMux I__793 (
            .O(N__4017),
            .I(N__4014));
    Span4Mux_s3_v I__792 (
            .O(N__4014),
            .I(N__4011));
    Span4Mux_v I__791 (
            .O(N__4011),
            .I(N__4008));
    Sp12to4 I__790 (
            .O(N__4008),
            .I(N__4005));
    Span12Mux_s10_h I__789 (
            .O(N__4005),
            .I(N__4002));
    Odrv12 I__788 (
            .O(N__4002),
            .I(lcol1_c));
    IoInMux I__787 (
            .O(N__3999),
            .I(N__3996));
    LocalMux I__786 (
            .O(N__3996),
            .I(N__3993));
    Span4Mux_s3_v I__785 (
            .O(N__3993),
            .I(N__3990));
    Sp12to4 I__784 (
            .O(N__3990),
            .I(N__3987));
    Span12Mux_h I__783 (
            .O(N__3987),
            .I(N__3984));
    Span12Mux_v I__782 (
            .O(N__3984),
            .I(N__3981));
    Odrv12 I__781 (
            .O(N__3981),
            .I(lcol2_c));
    IoInMux I__780 (
            .O(N__3978),
            .I(N__3975));
    LocalMux I__779 (
            .O(N__3975),
            .I(N__3972));
    Span4Mux_s3_v I__778 (
            .O(N__3972),
            .I(N__3969));
    Span4Mux_h I__777 (
            .O(N__3969),
            .I(N__3966));
    Span4Mux_v I__776 (
            .O(N__3966),
            .I(N__3963));
    Span4Mux_v I__775 (
            .O(N__3963),
            .I(N__3960));
    Span4Mux_v I__774 (
            .O(N__3960),
            .I(N__3957));
    Odrv4 I__773 (
            .O(N__3957),
            .I(lcol3_c));
    InMux I__772 (
            .O(N__3954),
            .I(N__3950));
    InMux I__771 (
            .O(N__3953),
            .I(N__3943));
    LocalMux I__770 (
            .O(N__3950),
            .I(N__3940));
    InMux I__769 (
            .O(N__3949),
            .I(N__3935));
    InMux I__768 (
            .O(N__3948),
            .I(N__3935));
    InMux I__767 (
            .O(N__3947),
            .I(N__3930));
    InMux I__766 (
            .O(N__3946),
            .I(N__3927));
    LocalMux I__765 (
            .O(N__3943),
            .I(N__3924));
    Span4Mux_v I__764 (
            .O(N__3940),
            .I(N__3919));
    LocalMux I__763 (
            .O(N__3935),
            .I(N__3919));
    CascadeMux I__762 (
            .O(N__3934),
            .I(N__3902));
    CascadeMux I__761 (
            .O(N__3933),
            .I(N__3895));
    LocalMux I__760 (
            .O(N__3930),
            .I(N__3890));
    LocalMux I__759 (
            .O(N__3927),
            .I(N__3890));
    Span4Mux_v I__758 (
            .O(N__3924),
            .I(N__3885));
    Span4Mux_v I__757 (
            .O(N__3919),
            .I(N__3885));
    InMux I__756 (
            .O(N__3918),
            .I(N__3882));
    InMux I__755 (
            .O(N__3917),
            .I(N__3875));
    InMux I__754 (
            .O(N__3916),
            .I(N__3875));
    InMux I__753 (
            .O(N__3915),
            .I(N__3875));
    InMux I__752 (
            .O(N__3914),
            .I(N__3872));
    InMux I__751 (
            .O(N__3913),
            .I(N__3861));
    InMux I__750 (
            .O(N__3912),
            .I(N__3861));
    InMux I__749 (
            .O(N__3911),
            .I(N__3861));
    InMux I__748 (
            .O(N__3910),
            .I(N__3861));
    InMux I__747 (
            .O(N__3909),
            .I(N__3861));
    InMux I__746 (
            .O(N__3908),
            .I(N__3856));
    InMux I__745 (
            .O(N__3907),
            .I(N__3856));
    InMux I__744 (
            .O(N__3906),
            .I(N__3849));
    InMux I__743 (
            .O(N__3905),
            .I(N__3849));
    InMux I__742 (
            .O(N__3902),
            .I(N__3849));
    InMux I__741 (
            .O(N__3901),
            .I(N__3844));
    InMux I__740 (
            .O(N__3900),
            .I(N__3844));
    InMux I__739 (
            .O(N__3899),
            .I(N__3837));
    InMux I__738 (
            .O(N__3898),
            .I(N__3837));
    InMux I__737 (
            .O(N__3895),
            .I(N__3837));
    Odrv4 I__736 (
            .O(N__3890),
            .I(colZ0Z_1));
    Odrv4 I__735 (
            .O(N__3885),
            .I(colZ0Z_1));
    LocalMux I__734 (
            .O(N__3882),
            .I(colZ0Z_1));
    LocalMux I__733 (
            .O(N__3875),
            .I(colZ0Z_1));
    LocalMux I__732 (
            .O(N__3872),
            .I(colZ0Z_1));
    LocalMux I__731 (
            .O(N__3861),
            .I(colZ0Z_1));
    LocalMux I__730 (
            .O(N__3856),
            .I(colZ0Z_1));
    LocalMux I__729 (
            .O(N__3849),
            .I(colZ0Z_1));
    LocalMux I__728 (
            .O(N__3844),
            .I(colZ0Z_1));
    LocalMux I__727 (
            .O(N__3837),
            .I(colZ0Z_1));
    CascadeMux I__726 (
            .O(N__3816),
            .I(N__3813));
    InMux I__725 (
            .O(N__3813),
            .I(N__3806));
    InMux I__724 (
            .O(N__3812),
            .I(N__3798));
    InMux I__723 (
            .O(N__3811),
            .I(N__3798));
    InMux I__722 (
            .O(N__3810),
            .I(N__3795));
    InMux I__721 (
            .O(N__3809),
            .I(N__3789));
    LocalMux I__720 (
            .O(N__3806),
            .I(N__3786));
    InMux I__719 (
            .O(N__3805),
            .I(N__3783));
    InMux I__718 (
            .O(N__3804),
            .I(N__3778));
    InMux I__717 (
            .O(N__3803),
            .I(N__3778));
    LocalMux I__716 (
            .O(N__3798),
            .I(N__3773));
    LocalMux I__715 (
            .O(N__3795),
            .I(N__3773));
    CascadeMux I__714 (
            .O(N__3794),
            .I(N__3770));
    CascadeMux I__713 (
            .O(N__3793),
            .I(N__3760));
    CascadeMux I__712 (
            .O(N__3792),
            .I(N__3757));
    LocalMux I__711 (
            .O(N__3789),
            .I(N__3744));
    Span4Mux_h I__710 (
            .O(N__3786),
            .I(N__3735));
    LocalMux I__709 (
            .O(N__3783),
            .I(N__3735));
    LocalMux I__708 (
            .O(N__3778),
            .I(N__3735));
    Span4Mux_v I__707 (
            .O(N__3773),
            .I(N__3735));
    InMux I__706 (
            .O(N__3770),
            .I(N__3732));
    InMux I__705 (
            .O(N__3769),
            .I(N__3729));
    InMux I__704 (
            .O(N__3768),
            .I(N__3722));
    InMux I__703 (
            .O(N__3767),
            .I(N__3722));
    InMux I__702 (
            .O(N__3766),
            .I(N__3722));
    InMux I__701 (
            .O(N__3765),
            .I(N__3719));
    InMux I__700 (
            .O(N__3764),
            .I(N__3714));
    InMux I__699 (
            .O(N__3763),
            .I(N__3714));
    InMux I__698 (
            .O(N__3760),
            .I(N__3709));
    InMux I__697 (
            .O(N__3757),
            .I(N__3709));
    InMux I__696 (
            .O(N__3756),
            .I(N__3704));
    InMux I__695 (
            .O(N__3755),
            .I(N__3704));
    InMux I__694 (
            .O(N__3754),
            .I(N__3697));
    InMux I__693 (
            .O(N__3753),
            .I(N__3697));
    InMux I__692 (
            .O(N__3752),
            .I(N__3697));
    InMux I__691 (
            .O(N__3751),
            .I(N__3692));
    InMux I__690 (
            .O(N__3750),
            .I(N__3692));
    InMux I__689 (
            .O(N__3749),
            .I(N__3685));
    InMux I__688 (
            .O(N__3748),
            .I(N__3685));
    InMux I__687 (
            .O(N__3747),
            .I(N__3685));
    Odrv4 I__686 (
            .O(N__3744),
            .I(colZ0Z_0));
    Odrv4 I__685 (
            .O(N__3735),
            .I(colZ0Z_0));
    LocalMux I__684 (
            .O(N__3732),
            .I(colZ0Z_0));
    LocalMux I__683 (
            .O(N__3729),
            .I(colZ0Z_0));
    LocalMux I__682 (
            .O(N__3722),
            .I(colZ0Z_0));
    LocalMux I__681 (
            .O(N__3719),
            .I(colZ0Z_0));
    LocalMux I__680 (
            .O(N__3714),
            .I(colZ0Z_0));
    LocalMux I__679 (
            .O(N__3709),
            .I(colZ0Z_0));
    LocalMux I__678 (
            .O(N__3704),
            .I(colZ0Z_0));
    LocalMux I__677 (
            .O(N__3697),
            .I(colZ0Z_0));
    LocalMux I__676 (
            .O(N__3692),
            .I(colZ0Z_0));
    LocalMux I__675 (
            .O(N__3685),
            .I(colZ0Z_0));
    IoInMux I__674 (
            .O(N__3660),
            .I(N__3657));
    LocalMux I__673 (
            .O(N__3657),
            .I(N__3654));
    IoSpan4Mux I__672 (
            .O(N__3654),
            .I(N__3651));
    Span4Mux_s1_v I__671 (
            .O(N__3651),
            .I(N__3648));
    Sp12to4 I__670 (
            .O(N__3648),
            .I(N__3645));
    Span12Mux_v I__669 (
            .O(N__3645),
            .I(N__3642));
    Span12Mux_h I__668 (
            .O(N__3642),
            .I(N__3639));
    Odrv12 I__667 (
            .O(N__3639),
            .I(lcol4_c));
    CEMux I__666 (
            .O(N__3636),
            .I(N__3633));
    LocalMux I__665 (
            .O(N__3633),
            .I(N__3630));
    Span4Mux_v I__664 (
            .O(N__3630),
            .I(N__3624));
    CEMux I__663 (
            .O(N__3629),
            .I(N__3621));
    CEMux I__662 (
            .O(N__3628),
            .I(N__3618));
    CEMux I__661 (
            .O(N__3627),
            .I(N__3615));
    Span4Mux_v I__660 (
            .O(N__3624),
            .I(N__3608));
    LocalMux I__659 (
            .O(N__3621),
            .I(N__3608));
    LocalMux I__658 (
            .O(N__3618),
            .I(N__3605));
    LocalMux I__657 (
            .O(N__3615),
            .I(N__3602));
    CEMux I__656 (
            .O(N__3614),
            .I(N__3599));
    CEMux I__655 (
            .O(N__3613),
            .I(N__3596));
    Span4Mux_v I__654 (
            .O(N__3608),
            .I(N__3593));
    Span4Mux_v I__653 (
            .O(N__3605),
            .I(N__3586));
    Span4Mux_v I__652 (
            .O(N__3602),
            .I(N__3586));
    LocalMux I__651 (
            .O(N__3599),
            .I(N__3586));
    LocalMux I__650 (
            .O(N__3596),
            .I(N__3577));
    Span4Mux_h I__649 (
            .O(N__3593),
            .I(N__3574));
    Span4Mux_v I__648 (
            .O(N__3586),
            .I(N__3571));
    InMux I__647 (
            .O(N__3585),
            .I(N__3564));
    InMux I__646 (
            .O(N__3584),
            .I(N__3564));
    InMux I__645 (
            .O(N__3583),
            .I(N__3564));
    InMux I__644 (
            .O(N__3582),
            .I(N__3559));
    InMux I__643 (
            .O(N__3581),
            .I(N__3559));
    InMux I__642 (
            .O(N__3580),
            .I(N__3556));
    Odrv12 I__641 (
            .O(N__3577),
            .I(clock_out_RNIR6ER_0));
    Odrv4 I__640 (
            .O(N__3574),
            .I(clock_out_RNIR6ER_0));
    Odrv4 I__639 (
            .O(N__3571),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__638 (
            .O(N__3564),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__637 (
            .O(N__3559),
            .I(clock_out_RNIR6ER_0));
    LocalMux I__636 (
            .O(N__3556),
            .I(clock_out_RNIR6ER_0));
    InMux I__635 (
            .O(N__3543),
            .I(N__3540));
    LocalMux I__634 (
            .O(N__3540),
            .I(N__3537));
    Span4Mux_v I__633 (
            .O(N__3537),
            .I(N__3534));
    Odrv4 I__632 (
            .O(N__3534),
            .I(delayConstant_fastZ0Z_2));
    InMux I__631 (
            .O(N__3531),
            .I(N__3528));
    LocalMux I__630 (
            .O(N__3528),
            .I(N__3525));
    Span4Mux_v I__629 (
            .O(N__3525),
            .I(N__3522));
    Odrv4 I__628 (
            .O(N__3522),
            .I(delayConstant_fastZ0Z_0));
    InMux I__627 (
            .O(N__3519),
            .I(N__3516));
    LocalMux I__626 (
            .O(N__3516),
            .I(\dig1.i2_mux ));
    InMux I__625 (
            .O(N__3513),
            .I(N__3510));
    LocalMux I__624 (
            .O(N__3510),
            .I(\dig1.m23_bm ));
    CascadeMux I__623 (
            .O(N__3507),
            .I(\dig1.m29_bm_cascade_ ));
    InMux I__622 (
            .O(N__3504),
            .I(N__3501));
    LocalMux I__621 (
            .O(N__3501),
            .I(\dig1.m23_am ));
    CascadeMux I__620 (
            .O(N__3498),
            .I(\dig1.m29_am_cascade_ ));
    InMux I__619 (
            .O(N__3495),
            .I(N__3492));
    LocalMux I__618 (
            .O(N__3492),
            .I(\dig1.m30_ns_1 ));
    CascadeMux I__617 (
            .O(N__3489),
            .I(N__3480));
    CascadeMux I__616 (
            .O(N__3488),
            .I(N__3477));
    CascadeMux I__615 (
            .O(N__3487),
            .I(N__3474));
    CascadeMux I__614 (
            .O(N__3486),
            .I(N__3471));
    InMux I__613 (
            .O(N__3485),
            .I(N__3462));
    InMux I__612 (
            .O(N__3484),
            .I(N__3459));
    InMux I__611 (
            .O(N__3483),
            .I(N__3449));
    InMux I__610 (
            .O(N__3480),
            .I(N__3449));
    InMux I__609 (
            .O(N__3477),
            .I(N__3449));
    InMux I__608 (
            .O(N__3474),
            .I(N__3449));
    InMux I__607 (
            .O(N__3471),
            .I(N__3444));
    InMux I__606 (
            .O(N__3470),
            .I(N__3444));
    CascadeMux I__605 (
            .O(N__3469),
            .I(N__3441));
    CascadeMux I__604 (
            .O(N__3468),
            .I(N__3437));
    CascadeMux I__603 (
            .O(N__3467),
            .I(N__3434));
    CascadeMux I__602 (
            .O(N__3466),
            .I(N__3431));
    CascadeMux I__601 (
            .O(N__3465),
            .I(N__3428));
    LocalMux I__600 (
            .O(N__3462),
            .I(N__3425));
    LocalMux I__599 (
            .O(N__3459),
            .I(N__3422));
    InMux I__598 (
            .O(N__3458),
            .I(N__3419));
    LocalMux I__597 (
            .O(N__3449),
            .I(N__3416));
    LocalMux I__596 (
            .O(N__3444),
            .I(N__3413));
    InMux I__595 (
            .O(N__3441),
            .I(N__3410));
    InMux I__594 (
            .O(N__3440),
            .I(N__3403));
    InMux I__593 (
            .O(N__3437),
            .I(N__3403));
    InMux I__592 (
            .O(N__3434),
            .I(N__3403));
    InMux I__591 (
            .O(N__3431),
            .I(N__3398));
    InMux I__590 (
            .O(N__3428),
            .I(N__3398));
    Odrv4 I__589 (
            .O(N__3425),
            .I(delayConstantZ0Z_0));
    Odrv12 I__588 (
            .O(N__3422),
            .I(delayConstantZ0Z_0));
    LocalMux I__587 (
            .O(N__3419),
            .I(delayConstantZ0Z_0));
    Odrv4 I__586 (
            .O(N__3416),
            .I(delayConstantZ0Z_0));
    Odrv4 I__585 (
            .O(N__3413),
            .I(delayConstantZ0Z_0));
    LocalMux I__584 (
            .O(N__3410),
            .I(delayConstantZ0Z_0));
    LocalMux I__583 (
            .O(N__3403),
            .I(delayConstantZ0Z_0));
    LocalMux I__582 (
            .O(N__3398),
            .I(delayConstantZ0Z_0));
    InMux I__581 (
            .O(N__3381),
            .I(N__3375));
    InMux I__580 (
            .O(N__3380),
            .I(N__3364));
    InMux I__579 (
            .O(N__3379),
            .I(N__3364));
    InMux I__578 (
            .O(N__3378),
            .I(N__3364));
    LocalMux I__577 (
            .O(N__3375),
            .I(N__3361));
    InMux I__576 (
            .O(N__3374),
            .I(N__3354));
    InMux I__575 (
            .O(N__3373),
            .I(N__3354));
    InMux I__574 (
            .O(N__3372),
            .I(N__3354));
    CascadeMux I__573 (
            .O(N__3371),
            .I(N__3351));
    LocalMux I__572 (
            .O(N__3364),
            .I(N__3348));
    Span4Mux_v I__571 (
            .O(N__3361),
            .I(N__3343));
    LocalMux I__570 (
            .O(N__3354),
            .I(N__3343));
    InMux I__569 (
            .O(N__3351),
            .I(N__3340));
    Odrv12 I__568 (
            .O(N__3348),
            .I(delayConstantZ0Z_2));
    Odrv4 I__567 (
            .O(N__3343),
            .I(delayConstantZ0Z_2));
    LocalMux I__566 (
            .O(N__3340),
            .I(delayConstantZ0Z_2));
    InMux I__565 (
            .O(N__3333),
            .I(N__3330));
    LocalMux I__564 (
            .O(N__3330),
            .I(N__3327));
    Odrv4 I__563 (
            .O(N__3327),
            .I(\dig1.leds_cnst_1 ));
    IoInMux I__562 (
            .O(N__3324),
            .I(N__3321));
    LocalMux I__561 (
            .O(N__3321),
            .I(N__3318));
    Span4Mux_s3_v I__560 (
            .O(N__3318),
            .I(N__3315));
    Span4Mux_v I__559 (
            .O(N__3315),
            .I(N__3312));
    Sp12to4 I__558 (
            .O(N__3312),
            .I(N__3309));
    Span12Mux_s10_h I__557 (
            .O(N__3309),
            .I(N__3306));
    Odrv12 I__556 (
            .O(N__3306),
            .I(leds_1_i_0_1));
    InMux I__555 (
            .O(N__3303),
            .I(N__3299));
    InMux I__554 (
            .O(N__3302),
            .I(N__3296));
    LocalMux I__553 (
            .O(N__3299),
            .I(un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2));
    LocalMux I__552 (
            .O(N__3296),
            .I(un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2));
    InMux I__551 (
            .O(N__3291),
            .I(N__3287));
    InMux I__550 (
            .O(N__3290),
            .I(N__3284));
    LocalMux I__549 (
            .O(N__3287),
            .I(un1_delayConstant_cry_3_0_c_RNITFZ0Z062));
    LocalMux I__548 (
            .O(N__3284),
            .I(un1_delayConstant_cry_3_0_c_RNITFZ0Z062));
    InMux I__547 (
            .O(N__3279),
            .I(N__3275));
    InMux I__546 (
            .O(N__3278),
            .I(N__3272));
    LocalMux I__545 (
            .O(N__3275),
            .I(un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2));
    LocalMux I__544 (
            .O(N__3272),
            .I(un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2));
    InMux I__543 (
            .O(N__3267),
            .I(N__3261));
    InMux I__542 (
            .O(N__3266),
            .I(N__3261));
    LocalMux I__541 (
            .O(N__3261),
            .I(un1_delayConstant_cry_1_0_c_RNIP5KDZ0Z2));
    CascadeMux I__540 (
            .O(N__3258),
            .I(\dig1.m8_am_cascade_ ));
    InMux I__539 (
            .O(N__3255),
            .I(N__3252));
    LocalMux I__538 (
            .O(N__3252),
            .I(\dig1.m8_bm ));
    CascadeMux I__537 (
            .O(N__3249),
            .I(\dig1.N_9_cascade_ ));
    CascadeMux I__536 (
            .O(N__3246),
            .I(clock_out_RNIR6ER_0_cascade_));
    CascadeMux I__535 (
            .O(N__3243),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4_cascade_ ));
    CascadeMux I__534 (
            .O(N__3240),
            .I(N__3235));
    CascadeMux I__533 (
            .O(N__3239),
            .I(N__3232));
    InMux I__532 (
            .O(N__3238),
            .I(N__3228));
    InMux I__531 (
            .O(N__3235),
            .I(N__3223));
    InMux I__530 (
            .O(N__3232),
            .I(N__3223));
    InMux I__529 (
            .O(N__3231),
            .I(N__3220));
    LocalMux I__528 (
            .O(N__3228),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4 ));
    LocalMux I__527 (
            .O(N__3223),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4 ));
    LocalMux I__526 (
            .O(N__3220),
            .I(\debounceconsolereset.counter_RNINST81Z0Z_4 ));
    IoInMux I__525 (
            .O(N__3213),
            .I(N__3210));
    LocalMux I__524 (
            .O(N__3210),
            .I(N__3207));
    Span4Mux_s0_v I__523 (
            .O(N__3207),
            .I(N__3204));
    Span4Mux_v I__522 (
            .O(N__3204),
            .I(N__3198));
    InMux I__521 (
            .O(N__3203),
            .I(N__3193));
    InMux I__520 (
            .O(N__3202),
            .I(N__3193));
    InMux I__519 (
            .O(N__3201),
            .I(N__3189));
    Span4Mux_v I__518 (
            .O(N__3198),
            .I(N__3183));
    LocalMux I__517 (
            .O(N__3193),
            .I(N__3183));
    InMux I__516 (
            .O(N__3192),
            .I(N__3180));
    LocalMux I__515 (
            .O(N__3189),
            .I(N__3177));
    InMux I__514 (
            .O(N__3188),
            .I(N__3174));
    Span4Mux_h I__513 (
            .O(N__3183),
            .I(N__3171));
    LocalMux I__512 (
            .O(N__3180),
            .I(N__3168));
    Span4Mux_v I__511 (
            .O(N__3177),
            .I(N__3165));
    LocalMux I__510 (
            .O(N__3174),
            .I(N__3162));
    Span4Mux_v I__509 (
            .O(N__3171),
            .I(N__3157));
    Span4Mux_h I__508 (
            .O(N__3168),
            .I(N__3157));
    Sp12to4 I__507 (
            .O(N__3165),
            .I(N__3154));
    Sp12to4 I__506 (
            .O(N__3162),
            .I(N__3151));
    Span4Mux_h I__505 (
            .O(N__3157),
            .I(N__3148));
    Span12Mux_h I__504 (
            .O(N__3154),
            .I(N__3145));
    Span12Mux_v I__503 (
            .O(N__3151),
            .I(N__3142));
    Sp12to4 I__502 (
            .O(N__3148),
            .I(N__3139));
    Span12Mux_v I__501 (
            .O(N__3145),
            .I(N__3136));
    Span12Mux_h I__500 (
            .O(N__3142),
            .I(N__3131));
    Span12Mux_v I__499 (
            .O(N__3139),
            .I(N__3131));
    Odrv12 I__498 (
            .O(N__3136),
            .I(masterreset_c));
    Odrv12 I__497 (
            .O(N__3131),
            .I(masterreset_c));
    InMux I__496 (
            .O(N__3126),
            .I(N__3117));
    InMux I__495 (
            .O(N__3125),
            .I(N__3117));
    InMux I__494 (
            .O(N__3124),
            .I(N__3117));
    LocalMux I__493 (
            .O(N__3117),
            .I(N__3113));
    CascadeMux I__492 (
            .O(N__3116),
            .I(N__3110));
    Span4Mux_v I__491 (
            .O(N__3113),
            .I(N__3106));
    InMux I__490 (
            .O(N__3110),
            .I(N__3101));
    InMux I__489 (
            .O(N__3109),
            .I(N__3101));
    Odrv4 I__488 (
            .O(N__3106),
            .I(slowclk));
    LocalMux I__487 (
            .O(N__3101),
            .I(slowclk));
    InMux I__486 (
            .O(N__3096),
            .I(N__3091));
    InMux I__485 (
            .O(N__3095),
            .I(N__3086));
    InMux I__484 (
            .O(N__3094),
            .I(N__3086));
    LocalMux I__483 (
            .O(N__3091),
            .I(debouncedn_counter_4));
    LocalMux I__482 (
            .O(N__3086),
            .I(debouncedn_counter_4));
    CascadeMux I__481 (
            .O(N__3081),
            .I(N__3078));
    InMux I__480 (
            .O(N__3078),
            .I(N__3073));
    InMux I__479 (
            .O(N__3077),
            .I(N__3068));
    InMux I__478 (
            .O(N__3076),
            .I(N__3068));
    LocalMux I__477 (
            .O(N__3073),
            .I(debouncedn_counter_1));
    LocalMux I__476 (
            .O(N__3068),
            .I(debouncedn_counter_1));
    CascadeMux I__475 (
            .O(N__3063),
            .I(N__3058));
    InMux I__474 (
            .O(N__3062),
            .I(N__3054));
    InMux I__473 (
            .O(N__3061),
            .I(N__3047));
    InMux I__472 (
            .O(N__3058),
            .I(N__3047));
    InMux I__471 (
            .O(N__3057),
            .I(N__3047));
    LocalMux I__470 (
            .O(N__3054),
            .I(debouncedn_counter_0));
    LocalMux I__469 (
            .O(N__3047),
            .I(debouncedn_counter_0));
    InMux I__468 (
            .O(N__3042),
            .I(N__3036));
    InMux I__467 (
            .O(N__3041),
            .I(N__3033));
    InMux I__466 (
            .O(N__3040),
            .I(N__3028));
    InMux I__465 (
            .O(N__3039),
            .I(N__3028));
    LocalMux I__464 (
            .O(N__3036),
            .I(N__3025));
    LocalMux I__463 (
            .O(N__3033),
            .I(debouncedn_counter_2));
    LocalMux I__462 (
            .O(N__3028),
            .I(debouncedn_counter_2));
    Odrv4 I__461 (
            .O(N__3025),
            .I(debouncedn_counter_2));
    InMux I__460 (
            .O(N__3018),
            .I(N__3015));
    LocalMux I__459 (
            .O(N__3015),
            .I(\debouncedn.out_cnvZ0Z_1 ));
    CascadeMux I__458 (
            .O(N__3012),
            .I(N__3008));
    CascadeMux I__457 (
            .O(N__3011),
            .I(N__3005));
    InMux I__456 (
            .O(N__3008),
            .I(N__3001));
    InMux I__455 (
            .O(N__3005),
            .I(N__2995));
    InMux I__454 (
            .O(N__3004),
            .I(N__2995));
    LocalMux I__453 (
            .O(N__3001),
            .I(N__2992));
    InMux I__452 (
            .O(N__3000),
            .I(N__2989));
    LocalMux I__451 (
            .O(N__2995),
            .I(debouncedn_counter_3));
    Odrv4 I__450 (
            .O(N__2992),
            .I(debouncedn_counter_3));
    LocalMux I__449 (
            .O(N__2989),
            .I(debouncedn_counter_3));
    InMux I__448 (
            .O(N__2982),
            .I(N__2979));
    LocalMux I__447 (
            .O(N__2979),
            .I(N__2976));
    Span4Mux_v I__446 (
            .O(N__2976),
            .I(N__2973));
    Sp12to4 I__445 (
            .O(N__2973),
            .I(N__2970));
    Span12Mux_h I__444 (
            .O(N__2970),
            .I(N__2967));
    Span12Mux_v I__443 (
            .O(N__2967),
            .I(N__2964));
    Odrv12 I__442 (
            .O(N__2964),
            .I(consolereset_c));
    InMux I__441 (
            .O(N__2961),
            .I(N__2958));
    LocalMux I__440 (
            .O(N__2958),
            .I(N__2955));
    Span4Mux_h I__439 (
            .O(N__2955),
            .I(N__2952));
    Sp12to4 I__438 (
            .O(N__2952),
            .I(N__2949));
    Span12Mux_v I__437 (
            .O(N__2949),
            .I(N__2946));
    Span12Mux_h I__436 (
            .O(N__2946),
            .I(N__2943));
    Odrv12 I__435 (
            .O(N__2943),
            .I(altreset_c));
    CascadeMux I__434 (
            .O(N__2940),
            .I(out_cnv_cascade_));
    CascadeMux I__433 (
            .O(N__2937),
            .I(col_1_1_cascade_));
    CascadeMux I__432 (
            .O(N__2934),
            .I(\dig1.m34_am_cascade_ ));
    InMux I__431 (
            .O(N__2931),
            .I(N__2928));
    LocalMux I__430 (
            .O(N__2928),
            .I(\dig1.m34_bm ));
    InMux I__429 (
            .O(N__2925),
            .I(\debounceconsolereset.un3_counter_cry_1 ));
    InMux I__428 (
            .O(N__2922),
            .I(\debounceconsolereset.un3_counter_cry_2 ));
    InMux I__427 (
            .O(N__2919),
            .I(\debounceconsolereset.un3_counter_cry_3 ));
    InMux I__426 (
            .O(N__2916),
            .I(N__2913));
    LocalMux I__425 (
            .O(N__2913),
            .I(\debounceconsolereset.un3_counter_cry_2_THRU_CO ));
    InMux I__424 (
            .O(N__2910),
            .I(N__2907));
    LocalMux I__423 (
            .O(N__2907),
            .I(\debounceconsolereset.un3_counter_cry_1_THRU_CO ));
    CascadeMux I__422 (
            .O(N__2904),
            .I(N__2900));
    CascadeMux I__421 (
            .O(N__2903),
            .I(N__2897));
    InMux I__420 (
            .O(N__2900),
            .I(N__2894));
    InMux I__419 (
            .O(N__2897),
            .I(N__2890));
    LocalMux I__418 (
            .O(N__2894),
            .I(N__2887));
    InMux I__417 (
            .O(N__2893),
            .I(N__2882));
    LocalMux I__416 (
            .O(N__2890),
            .I(N__2876));
    Span4Mux_h I__415 (
            .O(N__2887),
            .I(N__2873));
    InMux I__414 (
            .O(N__2886),
            .I(N__2870));
    InMux I__413 (
            .O(N__2885),
            .I(N__2867));
    LocalMux I__412 (
            .O(N__2882),
            .I(N__2864));
    InMux I__411 (
            .O(N__2881),
            .I(N__2859));
    InMux I__410 (
            .O(N__2880),
            .I(N__2859));
    InMux I__409 (
            .O(N__2879),
            .I(N__2856));
    Odrv4 I__408 (
            .O(N__2876),
            .I(delayConstantZ0Z_6));
    Odrv4 I__407 (
            .O(N__2873),
            .I(delayConstantZ0Z_6));
    LocalMux I__406 (
            .O(N__2870),
            .I(delayConstantZ0Z_6));
    LocalMux I__405 (
            .O(N__2867),
            .I(delayConstantZ0Z_6));
    Odrv4 I__404 (
            .O(N__2864),
            .I(delayConstantZ0Z_6));
    LocalMux I__403 (
            .O(N__2859),
            .I(delayConstantZ0Z_6));
    LocalMux I__402 (
            .O(N__2856),
            .I(delayConstantZ0Z_6));
    CascadeMux I__401 (
            .O(N__2841),
            .I(\dig2.m8_am_0_cascade_ ));
    InMux I__400 (
            .O(N__2838),
            .I(N__2835));
    LocalMux I__399 (
            .O(N__2835),
            .I(\dig2.N_9 ));
    CascadeMux I__398 (
            .O(N__2832),
            .I(slowclk_0_cascade_));
    CascadeMux I__397 (
            .O(N__2829),
            .I(N__2826));
    InMux I__396 (
            .O(N__2826),
            .I(N__2823));
    LocalMux I__395 (
            .O(N__2823),
            .I(slowclk_0));
    CascadeMux I__394 (
            .O(N__2820),
            .I(N__2811));
    CascadeMux I__393 (
            .O(N__2819),
            .I(N__2808));
    CascadeMux I__392 (
            .O(N__2818),
            .I(N__2803));
    CascadeMux I__391 (
            .O(N__2817),
            .I(N__2800));
    CascadeMux I__390 (
            .O(N__2816),
            .I(N__2797));
    CascadeMux I__389 (
            .O(N__2815),
            .I(N__2793));
    CascadeMux I__388 (
            .O(N__2814),
            .I(N__2790));
    InMux I__387 (
            .O(N__2811),
            .I(N__2784));
    InMux I__386 (
            .O(N__2808),
            .I(N__2784));
    CascadeMux I__385 (
            .O(N__2807),
            .I(N__2781));
    InMux I__384 (
            .O(N__2806),
            .I(N__2775));
    InMux I__383 (
            .O(N__2803),
            .I(N__2775));
    InMux I__382 (
            .O(N__2800),
            .I(N__2772));
    InMux I__381 (
            .O(N__2797),
            .I(N__2761));
    InMux I__380 (
            .O(N__2796),
            .I(N__2761));
    InMux I__379 (
            .O(N__2793),
            .I(N__2761));
    InMux I__378 (
            .O(N__2790),
            .I(N__2761));
    InMux I__377 (
            .O(N__2789),
            .I(N__2761));
    LocalMux I__376 (
            .O(N__2784),
            .I(N__2758));
    InMux I__375 (
            .O(N__2781),
            .I(N__2753));
    InMux I__374 (
            .O(N__2780),
            .I(N__2753));
    LocalMux I__373 (
            .O(N__2775),
            .I(delayConstantZ0Z_4));
    LocalMux I__372 (
            .O(N__2772),
            .I(delayConstantZ0Z_4));
    LocalMux I__371 (
            .O(N__2761),
            .I(delayConstantZ0Z_4));
    Odrv4 I__370 (
            .O(N__2758),
            .I(delayConstantZ0Z_4));
    LocalMux I__369 (
            .O(N__2753),
            .I(delayConstantZ0Z_4));
    CascadeMux I__368 (
            .O(N__2742),
            .I(N__2735));
    InMux I__367 (
            .O(N__2741),
            .I(N__2724));
    InMux I__366 (
            .O(N__2740),
            .I(N__2724));
    InMux I__365 (
            .O(N__2739),
            .I(N__2719));
    InMux I__364 (
            .O(N__2738),
            .I(N__2719));
    InMux I__363 (
            .O(N__2735),
            .I(N__2716));
    InMux I__362 (
            .O(N__2734),
            .I(N__2711));
    InMux I__361 (
            .O(N__2733),
            .I(N__2711));
    InMux I__360 (
            .O(N__2732),
            .I(N__2706));
    InMux I__359 (
            .O(N__2731),
            .I(N__2706));
    InMux I__358 (
            .O(N__2730),
            .I(N__2701));
    InMux I__357 (
            .O(N__2729),
            .I(N__2701));
    LocalMux I__356 (
            .O(N__2724),
            .I(N__2696));
    LocalMux I__355 (
            .O(N__2719),
            .I(N__2696));
    LocalMux I__354 (
            .O(N__2716),
            .I(delayConstantZ0Z_5));
    LocalMux I__353 (
            .O(N__2711),
            .I(delayConstantZ0Z_5));
    LocalMux I__352 (
            .O(N__2706),
            .I(delayConstantZ0Z_5));
    LocalMux I__351 (
            .O(N__2701),
            .I(delayConstantZ0Z_5));
    Odrv4 I__350 (
            .O(N__2696),
            .I(delayConstantZ0Z_5));
    InMux I__349 (
            .O(N__2685),
            .I(N__2682));
    LocalMux I__348 (
            .O(N__2682),
            .I(\dig2.m8_bm_0 ));
    InMux I__347 (
            .O(N__2679),
            .I(N__2675));
    InMux I__346 (
            .O(N__2678),
            .I(N__2672));
    LocalMux I__345 (
            .O(N__2675),
            .I(col_1_1));
    LocalMux I__344 (
            .O(N__2672),
            .I(col_1_1));
    InMux I__343 (
            .O(N__2667),
            .I(N__2664));
    LocalMux I__342 (
            .O(N__2664),
            .I(olddn_RNISQ7L1Z0Z_0));
    InMux I__341 (
            .O(N__2661),
            .I(un1_delayConstant_cry_1));
    CascadeMux I__340 (
            .O(N__2658),
            .I(N__2655));
    InMux I__339 (
            .O(N__2655),
            .I(N__2652));
    LocalMux I__338 (
            .O(N__2652),
            .I(olddn_RNISQ7L1Z0Z_3));
    InMux I__337 (
            .O(N__2649),
            .I(un1_delayConstant_cry_2));
    InMux I__336 (
            .O(N__2646),
            .I(N__2643));
    LocalMux I__335 (
            .O(N__2643),
            .I(olddn_RNISQ7L1Z0Z_1));
    InMux I__334 (
            .O(N__2640),
            .I(un1_delayConstant_cry_3));
    InMux I__333 (
            .O(N__2637),
            .I(N__2634));
    LocalMux I__332 (
            .O(N__2634),
            .I(olddn_RNISQ7LZ0Z1));
    InMux I__331 (
            .O(N__2631),
            .I(un1_delayConstant_cry_4));
    InMux I__330 (
            .O(N__2628),
            .I(N__2625));
    LocalMux I__329 (
            .O(N__2625),
            .I(olddn_RNISQ7L1Z0Z_4));
    InMux I__328 (
            .O(N__2622),
            .I(un1_delayConstant_cry_5));
    InMux I__327 (
            .O(N__2619),
            .I(un1_delayConstant_cry_6));
    InMux I__326 (
            .O(N__2616),
            .I(N__2608));
    InMux I__325 (
            .O(N__2615),
            .I(N__2605));
    CascadeMux I__324 (
            .O(N__2614),
            .I(N__2601));
    CascadeMux I__323 (
            .O(N__2613),
            .I(N__2598));
    CascadeMux I__322 (
            .O(N__2612),
            .I(N__2595));
    InMux I__321 (
            .O(N__2611),
            .I(N__2590));
    LocalMux I__320 (
            .O(N__2608),
            .I(N__2585));
    LocalMux I__319 (
            .O(N__2605),
            .I(N__2585));
    InMux I__318 (
            .O(N__2604),
            .I(N__2582));
    InMux I__317 (
            .O(N__2601),
            .I(N__2571));
    InMux I__316 (
            .O(N__2598),
            .I(N__2571));
    InMux I__315 (
            .O(N__2595),
            .I(N__2571));
    InMux I__314 (
            .O(N__2594),
            .I(N__2571));
    InMux I__313 (
            .O(N__2593),
            .I(N__2571));
    LocalMux I__312 (
            .O(N__2590),
            .I(delayConstant16_i));
    Odrv4 I__311 (
            .O(N__2585),
            .I(delayConstant16_i));
    LocalMux I__310 (
            .O(N__2582),
            .I(delayConstant16_i));
    LocalMux I__309 (
            .O(N__2571),
            .I(delayConstant16_i));
    CascadeMux I__308 (
            .O(N__2562),
            .I(N__2557));
    InMux I__307 (
            .O(N__2561),
            .I(N__2554));
    InMux I__306 (
            .O(N__2560),
            .I(N__2544));
    InMux I__305 (
            .O(N__2557),
            .I(N__2541));
    LocalMux I__304 (
            .O(N__2554),
            .I(N__2538));
    InMux I__303 (
            .O(N__2553),
            .I(N__2535));
    InMux I__302 (
            .O(N__2552),
            .I(N__2522));
    InMux I__301 (
            .O(N__2551),
            .I(N__2522));
    InMux I__300 (
            .O(N__2550),
            .I(N__2522));
    InMux I__299 (
            .O(N__2549),
            .I(N__2522));
    InMux I__298 (
            .O(N__2548),
            .I(N__2522));
    InMux I__297 (
            .O(N__2547),
            .I(N__2522));
    LocalMux I__296 (
            .O(N__2544),
            .I(olddn_RNI1J1RZ0));
    LocalMux I__295 (
            .O(N__2541),
            .I(olddn_RNI1J1RZ0));
    Odrv4 I__294 (
            .O(N__2538),
            .I(olddn_RNI1J1RZ0));
    LocalMux I__293 (
            .O(N__2535),
            .I(olddn_RNI1J1RZ0));
    LocalMux I__292 (
            .O(N__2522),
            .I(olddn_RNI1J1RZ0));
    CascadeMux I__291 (
            .O(N__2511),
            .I(delayConstant16_i_cascade_));
    InMux I__290 (
            .O(N__2508),
            .I(N__2505));
    LocalMux I__289 (
            .O(N__2505),
            .I(oldupZ0));
    InMux I__288 (
            .O(N__2502),
            .I(N__2499));
    LocalMux I__287 (
            .O(N__2499),
            .I(un1_delayConstant_cry_0_c_RNOZ0));
    CascadeMux I__286 (
            .O(N__2496),
            .I(N__2493));
    InMux I__285 (
            .O(N__2493),
            .I(N__2490));
    LocalMux I__284 (
            .O(N__2490),
            .I(olddn_RNISQ7L1Z0Z_2));
    InMux I__283 (
            .O(N__2487),
            .I(un1_delayConstant_cry_0));
    InMux I__282 (
            .O(N__2484),
            .I(N__2481));
    LocalMux I__281 (
            .O(N__2481),
            .I(\dig2.m23_am_0 ));
    InMux I__280 (
            .O(N__2478),
            .I(N__2475));
    LocalMux I__279 (
            .O(N__2475),
            .I(\dig2.m29_am_0 ));
    InMux I__278 (
            .O(N__2472),
            .I(N__2469));
    LocalMux I__277 (
            .O(N__2469),
            .I(\dig2.N_38 ));
    InMux I__276 (
            .O(N__2466),
            .I(N__2463));
    LocalMux I__275 (
            .O(N__2463),
            .I(\dig2.m23_bm_0 ));
    CascadeMux I__274 (
            .O(N__2460),
            .I(\dig2.m34_am_0_cascade_ ));
    InMux I__273 (
            .O(N__2457),
            .I(N__2454));
    LocalMux I__272 (
            .O(N__2454),
            .I(\dig2.m34_bm_0 ));
    InMux I__271 (
            .O(N__2451),
            .I(N__2448));
    LocalMux I__270 (
            .O(N__2448),
            .I(\dig2.N_35 ));
    CascadeMux I__269 (
            .O(N__2445),
            .I(\dig2.leds_cnst_2_cascade_ ));
    IoInMux I__268 (
            .O(N__2442),
            .I(N__2439));
    LocalMux I__267 (
            .O(N__2439),
            .I(N__2436));
    Span12Mux_s7_v I__266 (
            .O(N__2436),
            .I(N__2433));
    Span12Mux_v I__265 (
            .O(N__2433),
            .I(N__2430));
    Span12Mux_h I__264 (
            .O(N__2430),
            .I(N__2427));
    Odrv12 I__263 (
            .O(N__2427),
            .I(leds_1_i_2));
    InMux I__262 (
            .O(N__2424),
            .I(N__2421));
    LocalMux I__261 (
            .O(N__2421),
            .I(olddnZ0));
    InMux I__260 (
            .O(N__2418),
            .I(N__2412));
    InMux I__259 (
            .O(N__2417),
            .I(N__2412));
    LocalMux I__258 (
            .O(N__2412),
            .I(debounceddn));
    InMux I__257 (
            .O(N__2409),
            .I(N__2404));
    InMux I__256 (
            .O(N__2408),
            .I(N__2399));
    InMux I__255 (
            .O(N__2407),
            .I(N__2399));
    LocalMux I__254 (
            .O(N__2404),
            .I(\dig2.un1_leds114_0 ));
    LocalMux I__253 (
            .O(N__2399),
            .I(\dig2.un1_leds114_0 ));
    CascadeMux I__252 (
            .O(N__2394),
            .I(\dig2.i2_mux_cascade_ ));
    InMux I__251 (
            .O(N__2391),
            .I(N__2388));
    LocalMux I__250 (
            .O(N__2388),
            .I(\dig2.leds_cnst_1 ));
    CascadeMux I__249 (
            .O(N__2385),
            .I(\dig2.m29_bm_0_cascade_ ));
    InMux I__248 (
            .O(N__2382),
            .I(N__2379));
    LocalMux I__247 (
            .O(N__2379),
            .I(\dig2.m30_ns_1 ));
    IoInMux I__246 (
            .O(N__2376),
            .I(N__2373));
    LocalMux I__245 (
            .O(N__2373),
            .I(N__2370));
    IoSpan4Mux I__244 (
            .O(N__2370),
            .I(N__2367));
    Span4Mux_s2_v I__243 (
            .O(N__2367),
            .I(N__2364));
    Sp12to4 I__242 (
            .O(N__2364),
            .I(N__2361));
    Span12Mux_s10_v I__241 (
            .O(N__2361),
            .I(N__2358));
    Span12Mux_v I__240 (
            .O(N__2358),
            .I(N__2355));
    Span12Mux_h I__239 (
            .O(N__2355),
            .I(N__2352));
    Odrv12 I__238 (
            .O(N__2352),
            .I(\arse.divseven.io_0_D_IN_0 ));
    IoInMux I__237 (
            .O(N__2349),
            .I(N__2346));
    LocalMux I__236 (
            .O(N__2346),
            .I(N__2343));
    Span12Mux_s8_h I__235 (
            .O(N__2343),
            .I(N__2340));
    Odrv12 I__234 (
            .O(N__2340),
            .I(masterreset_c_i));
    IoInMux I__233 (
            .O(N__2337),
            .I(N__2334));
    LocalMux I__232 (
            .O(N__2334),
            .I(N__2331));
    IoSpan4Mux I__231 (
            .O(N__2331),
            .I(N__2328));
    Odrv4 I__230 (
            .O(N__2328),
            .I(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO));
    InMux I__229 (
            .O(N__2325),
            .I(N__2322));
    LocalMux I__228 (
            .O(N__2322),
            .I(N__2319));
    Span4Mux_v I__227 (
            .O(N__2319),
            .I(N__2316));
    Sp12to4 I__226 (
            .O(N__2316),
            .I(N__2313));
    Span12Mux_h I__225 (
            .O(N__2313),
            .I(N__2310));
    Span12Mux_v I__224 (
            .O(N__2310),
            .I(N__2307));
    Odrv12 I__223 (
            .O(N__2307),
            .I(deldn_c));
    IoInMux I__222 (
            .O(N__2304),
            .I(N__2301));
    LocalMux I__221 (
            .O(N__2301),
            .I(N__2298));
    Span4Mux_s0_v I__220 (
            .O(N__2298),
            .I(N__2295));
    Sp12to4 I__219 (
            .O(N__2295),
            .I(N__2292));
    Span12Mux_h I__218 (
            .O(N__2292),
            .I(N__2289));
    Span12Mux_v I__217 (
            .O(N__2289),
            .I(N__2286));
    Odrv12 I__216 (
            .O(N__2286),
            .I(leds_1_i_1));
    IoInMux I__215 (
            .O(N__2283),
            .I(N__2280));
    LocalMux I__214 (
            .O(N__2280),
            .I(N__2277));
    Span4Mux_s3_v I__213 (
            .O(N__2277),
            .I(N__2274));
    Span4Mux_v I__212 (
            .O(N__2274),
            .I(N__2271));
    Sp12to4 I__211 (
            .O(N__2271),
            .I(N__2268));
    Span12Mux_h I__210 (
            .O(N__2268),
            .I(N__2265));
    Span12Mux_v I__209 (
            .O(N__2265),
            .I(N__2262));
    Odrv12 I__208 (
            .O(N__2262),
            .I(leds_1_i_3));
    ClkMux I__207 (
            .O(N__2259),
            .I(N__2256));
    GlobalMux I__206 (
            .O(N__2256),
            .I(N__2253));
    gio2CtrlBuf I__205 (
            .O(N__2253),
            .I(\arse.un1_io_0_1_g ));
    IoInMux I__204 (
            .O(N__2250),
            .I(N__2247));
    LocalMux I__203 (
            .O(N__2247),
            .I(N__2244));
    Span4Mux_s1_v I__202 (
            .O(N__2244),
            .I(N__2241));
    Sp12to4 I__201 (
            .O(N__2241),
            .I(N__2238));
    Span12Mux_h I__200 (
            .O(N__2238),
            .I(N__2235));
    Span12Mux_v I__199 (
            .O(N__2235),
            .I(N__2232));
    Span12Mux_v I__198 (
            .O(N__2232),
            .I(N__2229));
    Odrv12 I__197 (
            .O(N__2229),
            .I(\top_pll_nrtthrth.PLLOUTCORE ));
    INV \INVarse.diveight.dout_0C  (
            .O(\INVarse.diveight.dout_0C_net ),
            .I(N__5397));
    INV \INVarse.apusynclatchedC  (
            .O(\INVarse.apusynclatchedC_net ),
            .I(N__2259));
    INV \INVarse.cpuclkresetC  (
            .O(\INVarse.cpuclkresetC_net ),
            .I(N__5393));
    INV \INVarse.divseven.dout_0C  (
            .O(\INVarse.divseven.dout_0C_net ),
            .I(N__5392));
    INV \INVarse.cpuresetcount_0C  (
            .O(\INVarse.cpuresetcount_0C_net ),
            .I(N__5389));
    INV \INVarse.cpuresetoutregC  (
            .O(\INVarse.cpuresetoutregC_net ),
            .I(N__5387));
    INV \INVarse.doingsevenC  (
            .O(\INVarse.doingsevenC_net ),
            .I(N__5388));
    defparam IN_MUX_bfv_21_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_11_0_));
    defparam IN_MUX_bfv_22_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_8_0_));
    defparam IN_MUX_bfv_23_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_10_0_));
    defparam IN_MUX_bfv_23_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_11_0_ (
            .carryinitin(\arses.un2_counter_cry_8 ),
            .carryinitout(bfn_23_11_0_));
    defparam IN_MUX_bfv_24_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_8_0_));
    ICE_GB \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5  (
            .USERSIGNALTOGLOBALBUFFER(N__2250),
            .GLOBALBUFFEROUTPUT(PLLOUTCORE_g));
    ICE_GB \arse.divseven.io_0_RNIIG08  (
            .USERSIGNALTOGLOBALBUFFER(N__2376),
            .GLOBALBUFFEROUTPUT(\arse.un1_io_0_1_g ));
    ICE_GB masterreset_ibuf_RNIKP26_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2349),
            .GLOBALBUFFEROUTPUT(masterreset_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam masterreset_ibuf_RNIKP26_LC_15_16_2.C_ON=1'b0;
    defparam masterreset_ibuf_RNIKP26_LC_15_16_2.SEQ_MODE=4'b0000;
    defparam masterreset_ibuf_RNIKP26_LC_15_16_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 masterreset_ibuf_RNIKP26_LC_15_16_2 (
            .in0(N__3188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(masterreset_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2.C_ON=1'b0;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2 (
            .in0(N__5316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.out_e_0_LC_19_10_0 .C_ON=1'b0;
    defparam \debouncedn.out_e_0_LC_19_10_0 .SEQ_MODE=4'b1000;
    defparam \debouncedn.out_e_0_LC_19_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \debouncedn.out_e_0_LC_19_10_0  (
            .in0(N__2325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debounceddn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5293),
            .ce(N__5237),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_1_LC_19_12_0 .C_ON=1'b0;
    defparam \dig2.leds_1_i_1_LC_19_12_0 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_1_LC_19_12_0 .LUT_INIT=16'b0101010100000011;
    LogicCell40 \dig2.leds_1_i_1_LC_19_12_0  (
            .in0(N__2391),
            .in1(N__3953),
            .in2(N__3816),
            .in3(N__2409),
            .lcout(leds_1_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5297),
            .ce(N__3629),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_3_LC_19_13_0 .C_ON=1'b0;
    defparam \dig2.leds_1_i_3_LC_19_13_0 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_3_LC_19_13_0 .LUT_INIT=16'b1000000010001100;
    LogicCell40 \dig2.leds_1_i_3_LC_19_13_0  (
            .in0(N__2472),
            .in1(N__2408),
            .in2(N__5076),
            .in3(N__2451),
            .lcout(leds_1_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5300),
            .ce(N__3636),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m30_ns_LC_19_13_5 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m30_ns_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m30_ns_LC_19_13_5 .LUT_INIT=16'b0000101011111100;
    LogicCell40 \dig2.leds_cnst_3_1__m30_ns_LC_19_13_5  (
            .in0(N__2484),
            .in1(N__2478),
            .in2(N__2904),
            .in3(N__2382),
            .lcout(),
            .ltout(\dig2.leds_cnst_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_2_LC_19_13_6 .C_ON=1'b0;
    defparam \dig2.leds_1_i_2_LC_19_13_6 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_2_LC_19_13_6 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \dig2.leds_1_i_2_LC_19_13_6  (
            .in0(_gnd_net_),
            .in1(N__2407),
            .in2(N__2445),
            .in3(N__3809),
            .lcout(leds_1_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5300),
            .ce(N__3636),
            .sr(_gnd_net_));
    defparam olddn_LC_20_10_0.C_ON=1'b0;
    defparam olddn_LC_20_10_0.SEQ_MODE=4'b1000;
    defparam olddn_LC_20_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 olddn_LC_20_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2418),
            .lcout(olddnZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5294),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNI1J1R_LC_20_10_2.C_ON=1'b0;
    defparam olddn_RNI1J1R_LC_20_10_2.SEQ_MODE=4'b0000;
    defparam olddn_RNI1J1R_LC_20_10_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 olddn_RNI1J1R_LC_20_10_2 (
            .in0(_gnd_net_),
            .in1(N__2424),
            .in2(_gnd_net_),
            .in3(N__2417),
            .lcout(olddn_RNI1J1RZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNISQ7L1_3_LC_20_11_1.C_ON=1'b0;
    defparam olddn_RNISQ7L1_3_LC_20_11_1.SEQ_MODE=4'b0000;
    defparam olddn_RNISQ7L1_3_LC_20_11_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNISQ7L1_3_LC_20_11_1 (
            .in0(_gnd_net_),
            .in1(N__2604),
            .in2(_gnd_net_),
            .in3(N__2553),
            .lcout(olddn_RNISQ7L1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.un1_leds114_LC_20_12_2 .C_ON=1'b0;
    defparam \dig2.un1_leds114_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \dig2.un1_leds114_LC_20_12_2 .LUT_INIT=16'b1011110111111111;
    LogicCell40 \dig2.un1_leds114_LC_20_12_2  (
            .in0(N__2886),
            .in1(N__2806),
            .in2(N__5070),
            .in3(N__2734),
            .lcout(\dig2.un1_leds114_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m11_LC_20_12_3 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m11_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m11_LC_20_12_3 .LUT_INIT=16'b0001110011100011;
    LogicCell40 \dig2.leds_cnst_3_1__m11_LC_20_12_3  (
            .in0(N__2733),
            .in1(N__3918),
            .in2(N__2818),
            .in3(N__3769),
            .lcout(),
            .ltout(\dig2.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m13_LC_20_12_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m13_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m13_LC_20_12_4 .LUT_INIT=16'b1010001011110111;
    LogicCell40 \dig2.leds_cnst_3_1__m13_LC_20_12_4  (
            .in0(N__5056),
            .in1(N__2885),
            .in2(N__2394),
            .in3(N__2838),
            .lcout(\dig2.leds_cnst_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m29_bm_LC_20_13_0 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m29_bm_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m29_bm_LC_20_13_0 .LUT_INIT=16'b0110101001011101;
    LogicCell40 \dig2.leds_cnst_3_1__m29_bm_LC_20_13_0  (
            .in0(N__3766),
            .in1(N__2731),
            .in2(N__2814),
            .in3(N__3910),
            .lcout(),
            .ltout(\dig2.m29_bm_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m30_ns_1_LC_20_13_1 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m30_ns_1_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m30_ns_1_LC_20_13_1 .LUT_INIT=16'b0001100100111011;
    LogicCell40 \dig2.leds_cnst_3_1__m30_ns_1_LC_20_13_1  (
            .in0(N__2880),
            .in1(N__5071),
            .in2(N__2385),
            .in3(N__2466),
            .lcout(\dig2.m30_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m23_am_LC_20_13_3 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m23_am_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m23_am_LC_20_13_3 .LUT_INIT=16'b1111011110101101;
    LogicCell40 \dig2.leds_cnst_3_1__m23_am_LC_20_13_3  (
            .in0(N__3911),
            .in1(N__2730),
            .in2(N__3793),
            .in3(N__2796),
            .lcout(\dig2.m23_am_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m29_am_LC_20_13_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m29_am_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m29_am_LC_20_13_4 .LUT_INIT=16'b0101011101010101;
    LogicCell40 \dig2.leds_cnst_3_1__m29_am_LC_20_13_4  (
            .in0(N__3767),
            .in1(N__2732),
            .in2(N__2815),
            .in3(N__3912),
            .lcout(\dig2.m29_am_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m37_LC_20_13_6 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m37_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m37_LC_20_13_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \dig2.leds_cnst_3_1__m37_LC_20_13_6  (
            .in0(N__3768),
            .in1(N__3913),
            .in2(N__2816),
            .in3(N__2881),
            .lcout(\dig2.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m23_bm_LC_20_13_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m23_bm_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m23_bm_LC_20_13_7 .LUT_INIT=16'b0010011100000110;
    LogicCell40 \dig2.leds_cnst_3_1__m23_bm_LC_20_13_7  (
            .in0(N__3909),
            .in1(N__2729),
            .in2(N__3792),
            .in3(N__2789),
            .lcout(\dig2.m23_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m34_bm_LC_20_14_1 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m34_bm_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m34_bm_LC_20_14_1 .LUT_INIT=16'b0101000100110111;
    LogicCell40 \dig2.leds_cnst_3_1__m34_bm_LC_20_14_1  (
            .in0(N__2740),
            .in1(N__3914),
            .in2(N__2819),
            .in3(N__3765),
            .lcout(\dig2.m34_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m34_am_LC_20_14_5 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m34_am_LC_20_14_5 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m34_am_LC_20_14_5 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \dig2.leds_cnst_3_1__m34_am_LC_20_14_5  (
            .in0(N__2741),
            .in1(_gnd_net_),
            .in2(N__2820),
            .in3(N__2678),
            .lcout(),
            .ltout(\dig2.m34_am_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m34_ns_LC_20_14_6 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m34_ns_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m34_ns_LC_20_14_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \dig2.leds_cnst_3_1__m34_ns_LC_20_14_6  (
            .in0(_gnd_net_),
            .in1(N__2893),
            .in2(N__2460),
            .in3(N__2457),
            .lcout(\dig2.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_fast_0_LC_21_9_1.C_ON=1'b0;
    defparam delayConstant_fast_0_LC_21_9_1.SEQ_MODE=4'b1000;
    defparam delayConstant_fast_0_LC_21_9_1.LUT_INIT=16'b0101010110011001;
    LogicCell40 delayConstant_fast_0_LC_21_9_1 (
            .in0(N__3484),
            .in1(N__2611),
            .in2(_gnd_net_),
            .in3(N__2560),
            .lcout(delayConstant_fastZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5295),
            .ce(),
            .sr(N__4444));
    defparam \arses.counter_1_LC_21_9_7 .C_ON=1'b0;
    defparam \arses.counter_1_LC_21_9_7 .SEQ_MODE=4'b1001;
    defparam \arses.counter_1_LC_21_9_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \arses.counter_1_LC_21_9_7  (
            .in0(N__4132),
            .in1(N__4167),
            .in2(_gnd_net_),
            .in3(N__4557),
            .lcout(\arses.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5295),
            .ce(),
            .sr(N__4444));
    defparam olddn_RNISQ7L1_0_LC_21_10_0.C_ON=1'b0;
    defparam olddn_RNISQ7L1_0_LC_21_10_0.SEQ_MODE=4'b0000;
    defparam olddn_RNISQ7L1_0_LC_21_10_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNISQ7L1_0_LC_21_10_0 (
            .in0(_gnd_net_),
            .in1(N__2594),
            .in2(_gnd_net_),
            .in3(N__2549),
            .lcout(olddn_RNISQ7L1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam oldup_RNIR76Q_LC_21_10_1.C_ON=1'b0;
    defparam oldup_RNIR76Q_LC_21_10_1.SEQ_MODE=4'b0000;
    defparam oldup_RNIR76Q_LC_21_10_1.LUT_INIT=16'b1111111101110111;
    LogicCell40 oldup_RNIR76Q_LC_21_10_1 (
            .in0(N__3201),
            .in1(N__2508),
            .in2(_gnd_net_),
            .in3(N__5327),
            .lcout(delayConstant16_i),
            .ltout(delayConstant16_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_0_c_RNO_LC_21_10_2.C_ON=1'b0;
    defparam un1_delayConstant_cry_0_c_RNO_LC_21_10_2.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_0_c_RNO_LC_21_10_2.LUT_INIT=16'b1111111100001111;
    LogicCell40 un1_delayConstant_cry_0_c_RNO_LC_21_10_2 (
            .in0(N__3485),
            .in1(_gnd_net_),
            .in2(N__2511),
            .in3(N__2547),
            .lcout(un1_delayConstant_cry_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNISQ7L1_LC_21_10_3.C_ON=1'b0;
    defparam olddn_RNISQ7L1_LC_21_10_3.SEQ_MODE=4'b0000;
    defparam olddn_RNISQ7L1_LC_21_10_3.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNISQ7L1_LC_21_10_3 (
            .in0(N__2551),
            .in1(_gnd_net_),
            .in2(N__2613),
            .in3(_gnd_net_),
            .lcout(olddn_RNISQ7LZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam oldup_LC_21_10_4.C_ON=1'b0;
    defparam oldup_LC_21_10_4.SEQ_MODE=4'b1000;
    defparam oldup_LC_21_10_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 oldup_LC_21_10_4 (
            .in0(N__5328),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(oldupZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5298),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNISQ7L1_1_LC_21_10_5.C_ON=1'b0;
    defparam olddn_RNISQ7L1_1_LC_21_10_5.SEQ_MODE=4'b0000;
    defparam olddn_RNISQ7L1_1_LC_21_10_5.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNISQ7L1_1_LC_21_10_5 (
            .in0(N__2550),
            .in1(_gnd_net_),
            .in2(N__2612),
            .in3(_gnd_net_),
            .lcout(olddn_RNISQ7L1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNISQ7L1_2_LC_21_10_6.C_ON=1'b0;
    defparam olddn_RNISQ7L1_2_LC_21_10_6.SEQ_MODE=4'b0000;
    defparam olddn_RNISQ7L1_2_LC_21_10_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNISQ7L1_2_LC_21_10_6 (
            .in0(_gnd_net_),
            .in1(N__2593),
            .in2(_gnd_net_),
            .in3(N__2548),
            .lcout(olddn_RNISQ7L1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNISQ7L1_4_LC_21_10_7.C_ON=1'b0;
    defparam olddn_RNISQ7L1_4_LC_21_10_7.SEQ_MODE=4'b0000;
    defparam olddn_RNISQ7L1_4_LC_21_10_7.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNISQ7L1_4_LC_21_10_7 (
            .in0(N__2552),
            .in1(_gnd_net_),
            .in2(N__2614),
            .in3(_gnd_net_),
            .lcout(olddn_RNISQ7L1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_0_c_LC_21_11_0.C_ON=1'b1;
    defparam un1_delayConstant_cry_0_c_LC_21_11_0.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_0_c_LC_21_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_delayConstant_cry_0_c_LC_21_11_0 (
            .in0(_gnd_net_),
            .in1(N__2502),
            .in2(N__3469),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_11_0_),
            .carryout(un1_delayConstant_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_1_LC_21_11_1.C_ON=1'b1;
    defparam delayConstant_1_LC_21_11_1.SEQ_MODE=4'b1000;
    defparam delayConstant_1_LC_21_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_1_LC_21_11_1 (
            .in0(_gnd_net_),
            .in1(N__4979),
            .in2(N__2496),
            .in3(N__2487),
            .lcout(delayConstantZ0Z_1),
            .ltout(),
            .carryin(un1_delayConstant_cry_0),
            .carryout(un1_delayConstant_cry_1),
            .clk(N__5301),
            .ce(),
            .sr(N__4442));
    defparam un1_delayConstant_cry_1_0_c_RNIP5KD2_LC_21_11_2.C_ON=1'b1;
    defparam un1_delayConstant_cry_1_0_c_RNIP5KD2_LC_21_11_2.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_1_0_c_RNIP5KD2_LC_21_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_delayConstant_cry_1_0_c_RNIP5KD2_LC_21_11_2 (
            .in0(_gnd_net_),
            .in1(N__2667),
            .in2(N__3371),
            .in3(N__2661),
            .lcout(un1_delayConstant_cry_1_0_c_RNIP5KDZ0Z2),
            .ltout(),
            .carryin(un1_delayConstant_cry_1),
            .carryout(un1_delayConstant_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_3_LC_21_11_3.C_ON=1'b1;
    defparam delayConstant_3_LC_21_11_3.SEQ_MODE=4'b1000;
    defparam delayConstant_3_LC_21_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_3_LC_21_11_3 (
            .in0(_gnd_net_),
            .in1(N__4795),
            .in2(N__2658),
            .in3(N__2649),
            .lcout(delayConstantZ0Z_3),
            .ltout(),
            .carryin(un1_delayConstant_cry_2),
            .carryout(un1_delayConstant_cry_3),
            .clk(N__5301),
            .ce(),
            .sr(N__4442));
    defparam un1_delayConstant_cry_3_0_c_RNITF062_LC_21_11_4.C_ON=1'b1;
    defparam un1_delayConstant_cry_3_0_c_RNITF062_LC_21_11_4.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_3_0_c_RNITF062_LC_21_11_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_delayConstant_cry_3_0_c_RNITF062_LC_21_11_4 (
            .in0(_gnd_net_),
            .in1(N__2646),
            .in2(N__2817),
            .in3(N__2640),
            .lcout(un1_delayConstant_cry_3_0_c_RNITFZ0Z062),
            .ltout(),
            .carryin(un1_delayConstant_cry_3),
            .carryout(un1_delayConstant_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_4_0_c_RNIVK6A2_LC_21_11_5.C_ON=1'b1;
    defparam un1_delayConstant_cry_4_0_c_RNIVK6A2_LC_21_11_5.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_4_0_c_RNIVK6A2_LC_21_11_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_delayConstant_cry_4_0_c_RNIVK6A2_LC_21_11_5 (
            .in0(_gnd_net_),
            .in1(N__2637),
            .in2(N__2742),
            .in3(N__2631),
            .lcout(un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2),
            .ltout(),
            .carryin(un1_delayConstant_cry_4),
            .carryout(un1_delayConstant_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_5_0_c_RNI1QCE2_LC_21_11_6.C_ON=1'b1;
    defparam un1_delayConstant_cry_5_0_c_RNI1QCE2_LC_21_11_6.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_5_0_c_RNI1QCE2_LC_21_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_delayConstant_cry_5_0_c_RNI1QCE2_LC_21_11_6 (
            .in0(_gnd_net_),
            .in1(N__2628),
            .in2(N__2903),
            .in3(N__2622),
            .lcout(un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2),
            .ltout(),
            .carryin(un1_delayConstant_cry_5),
            .carryout(un1_delayConstant_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_7_LC_21_11_7.C_ON=1'b0;
    defparam delayConstant_7_LC_21_11_7.SEQ_MODE=4'b1000;
    defparam delayConstant_7_LC_21_11_7.LUT_INIT=16'b1001010101101010;
    LogicCell40 delayConstant_7_LC_21_11_7 (
            .in0(N__5060),
            .in1(N__2616),
            .in2(N__2562),
            .in3(N__2619),
            .lcout(delayConstantZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5301),
            .ce(),
            .sr(N__4442));
    defparam delayConstant_0_LC_21_12_1.C_ON=1'b0;
    defparam delayConstant_0_LC_21_12_1.SEQ_MODE=4'b1000;
    defparam delayConstant_0_LC_21_12_1.LUT_INIT=16'b0101010110011001;
    LogicCell40 delayConstant_0_LC_21_12_1 (
            .in0(N__3458),
            .in1(N__2615),
            .in2(_gnd_net_),
            .in3(N__2561),
            .lcout(delayConstantZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5303),
            .ce(),
            .sr(N__4441));
    defparam delayConstant_5_LC_21_12_4.C_ON=1'b0;
    defparam delayConstant_5_LC_21_12_4.SEQ_MODE=4'b1001;
    defparam delayConstant_5_LC_21_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_5_LC_21_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3278),
            .lcout(delayConstantZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5303),
            .ce(),
            .sr(N__4441));
    defparam delayConstant_4_LC_21_12_5.C_ON=1'b0;
    defparam delayConstant_4_LC_21_12_5.SEQ_MODE=4'b1000;
    defparam delayConstant_4_LC_21_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_4_LC_21_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3290),
            .lcout(delayConstantZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5303),
            .ce(),
            .sr(N__4441));
    defparam delayConstant_6_LC_21_12_7.C_ON=1'b0;
    defparam delayConstant_6_LC_21_12_7.SEQ_MODE=4'b1000;
    defparam delayConstant_6_LC_21_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_6_LC_21_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3302),
            .lcout(delayConstantZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5303),
            .ce(),
            .sr(N__4441));
    defparam \dig2.leds_cnst_3_1__m8_am_LC_21_13_0 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m8_am_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m8_am_LC_21_13_0 .LUT_INIT=16'b1101000001111010;
    LogicCell40 \dig2.leds_cnst_3_1__m8_am_LC_21_13_0  (
            .in0(N__2739),
            .in1(N__3898),
            .in2(N__2807),
            .in3(N__3748),
            .lcout(),
            .ltout(\dig2.m8_am_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m8_ns_LC_21_13_1 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m8_ns_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m8_ns_LC_21_13_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \dig2.leds_cnst_3_1__m8_ns_LC_21_13_1  (
            .in0(N__2879),
            .in1(_gnd_net_),
            .in2(N__2841),
            .in3(N__2685),
            .lcout(\dig2.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_LC_21_13_3 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_LC_21_13_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \arses.clock_out_RNIR6ER_LC_21_13_3  (
            .in0(N__3192),
            .in1(N__3124),
            .in2(_gnd_net_),
            .in3(N__4555),
            .lcout(slowclk_0),
            .ltout(slowclk_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam col_0_LC_21_13_4.C_ON=1'b0;
    defparam col_0_LC_21_13_4.SEQ_MODE=4'b1000;
    defparam col_0_LC_21_13_4.LUT_INIT=16'b1111010100001010;
    LogicCell40 col_0_LC_21_13_4 (
            .in0(N__3125),
            .in1(_gnd_net_),
            .in2(N__2832),
            .in3(N__3749),
            .lcout(colZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam col_1_LC_21_13_5.C_ON=1'b0;
    defparam col_1_LC_21_13_5.SEQ_MODE=4'b1000;
    defparam col_1_LC_21_13_5.LUT_INIT=16'b1010110010101010;
    LogicCell40 col_1_LC_21_13_5 (
            .in0(N__3899),
            .in1(N__2679),
            .in2(N__2829),
            .in3(N__3126),
            .lcout(colZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m8_bm_LC_21_13_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m8_bm_LC_21_13_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m8_bm_LC_21_13_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \dig2.leds_cnst_3_1__m8_bm_LC_21_13_7  (
            .in0(N__3747),
            .in1(N__2780),
            .in2(N__3933),
            .in3(N__2738),
            .lcout(\dig2.m8_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m34_bm_LC_21_14_2 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m34_bm_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m34_bm_LC_21_14_2 .LUT_INIT=16'b0101000100110111;
    LogicCell40 \dig1.leds_cnst_3_1__m34_bm_LC_21_14_2  (
            .in0(N__4993),
            .in1(N__3908),
            .in2(N__3486),
            .in3(N__3756),
            .lcout(\dig1.m34_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m11x_i_o2_LC_21_14_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m11x_i_o2_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m11x_i_o2_LC_21_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dig1.leds_cnst_3_1__m11x_i_o2_LC_21_14_4  (
            .in0(_gnd_net_),
            .in1(N__3907),
            .in2(_gnd_net_),
            .in3(N__3755),
            .lcout(col_1_1),
            .ltout(col_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m34_am_LC_21_14_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m34_am_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m34_am_LC_21_14_5 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \dig1.leds_cnst_3_1__m34_am_LC_21_14_5  (
            .in0(_gnd_net_),
            .in1(N__3470),
            .in2(N__2937),
            .in3(N__4994),
            .lcout(),
            .ltout(\dig1.m34_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m34_ns_LC_21_14_6 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m34_ns_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m34_ns_LC_21_14_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \dig1.leds_cnst_3_1__m34_ns_LC_21_14_6  (
            .in0(_gnd_net_),
            .in1(N__3381),
            .in2(N__2934),
            .in3(N__2931),
            .lcout(\dig1.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_22_8_0 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_22_8_0 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_22_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_1_c_LC_22_8_0  (
            .in0(_gnd_net_),
            .in1(N__3062),
            .in2(N__3081),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_8_0_),
            .carryout(\debounceconsolereset.un3_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_22_8_1 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_22_8_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_22_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_22_8_1  (
            .in0(_gnd_net_),
            .in1(N__3039),
            .in2(_gnd_net_),
            .in3(N__2925),
            .lcout(\debounceconsolereset.un3_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_1 ),
            .carryout(\debounceconsolereset.un3_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_22_8_2 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_22_8_2 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_22_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_22_8_2  (
            .in0(_gnd_net_),
            .in1(N__3004),
            .in2(_gnd_net_),
            .in3(N__2922),
            .lcout(\debounceconsolereset.un3_counter_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_2 ),
            .carryout(\debounceconsolereset.un3_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_4_LC_22_8_3 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_4_LC_22_8_3 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_4_LC_22_8_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \debounceconsolereset.counter_4_LC_22_8_3  (
            .in0(N__3096),
            .in1(N__3583),
            .in2(N__3239),
            .in3(N__2919),
            .lcout(debouncedn_counter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5296),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_3_LC_22_8_5 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_3_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_3_LC_22_8_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \debounceconsolereset.counter_3_LC_22_8_5  (
            .in0(N__2916),
            .in1(N__3585),
            .in2(N__3011),
            .in3(N__3238),
            .lcout(debouncedn_counter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5296),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_2_LC_22_8_7 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_2_LC_22_8_7 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_2_LC_22_8_7 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \debounceconsolereset.counter_2_LC_22_8_7  (
            .in0(N__2910),
            .in1(N__3584),
            .in2(N__3240),
            .in3(N__3040),
            .lcout(debouncedn_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5296),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_0_LC_22_9_0 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_0_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_0_LC_22_9_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \arses.clock_out_RNIR6ER_0_LC_22_9_0  (
            .in0(N__3203),
            .in1(N__3109),
            .in2(_gnd_net_),
            .in3(N__4500),
            .lcout(clock_out_RNIR6ER_0),
            .ltout(clock_out_RNIR6ER_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNINST81_4_LC_22_9_1 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_RNINST81_4_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNINST81_4_LC_22_9_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \debounceconsolereset.counter_RNINST81_4_LC_22_9_1  (
            .in0(N__3095),
            .in1(N__3000),
            .in2(N__3246),
            .in3(N__3041),
            .lcout(\debounceconsolereset.counter_RNINST81Z0Z_4 ),
            .ltout(\debounceconsolereset.counter_RNINST81Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_0_LC_22_9_2 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_0_LC_22_9_2 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_0_LC_22_9_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \debounceconsolereset.counter_0_LC_22_9_2  (
            .in0(N__3061),
            .in1(_gnd_net_),
            .in2(N__3243),
            .in3(N__3581),
            .lcout(debouncedn_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5299),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_1_LC_22_9_4 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_1_LC_22_9_4 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_1_LC_22_9_4 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \debounceconsolereset.counter_1_LC_22_9_4  (
            .in0(N__3077),
            .in1(N__3231),
            .in2(N__3063),
            .in3(N__3582),
            .lcout(debouncedn_counter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5299),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_LC_22_9_5 .C_ON=1'b0;
    defparam \arses.clock_out_LC_22_9_5 .SEQ_MODE=4'b1000;
    defparam \arses.clock_out_LC_22_9_5 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \arses.clock_out_LC_22_9_5  (
            .in0(N__4501),
            .in1(_gnd_net_),
            .in2(N__3116),
            .in3(N__3202),
            .lcout(slowclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5299),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.out_cnv_1_LC_22_9_7 .C_ON=1'b0;
    defparam \debouncedn.out_cnv_1_LC_22_9_7 .SEQ_MODE=4'b0000;
    defparam \debouncedn.out_cnv_1_LC_22_9_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \debouncedn.out_cnv_1_LC_22_9_7  (
            .in0(N__3094),
            .in1(N__3076),
            .in2(_gnd_net_),
            .in3(N__3057),
            .lcout(\debouncedn.out_cnvZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI1L5_2_LC_22_10_2 .C_ON=1'b0;
    defparam \arses.counter_RNI1L5_2_LC_22_10_2 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI1L5_2_LC_22_10_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \arses.counter_RNI1L5_2_LC_22_10_2  (
            .in0(N__4343),
            .in1(N__4112),
            .in2(_gnd_net_),
            .in3(N__4161),
            .lcout(\arses.un1_counterlto4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.out_cnv_LC_22_10_4 .C_ON=1'b0;
    defparam \debouncedn.out_cnv_LC_22_10_4 .SEQ_MODE=4'b0000;
    defparam \debouncedn.out_cnv_LC_22_10_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \debouncedn.out_cnv_LC_22_10_4  (
            .in0(N__3042),
            .in1(N__3018),
            .in2(N__3012),
            .in3(N__3580),
            .lcout(out_cnv),
            .ltout(out_cnv_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_LC_22_10_5 .C_ON=1'b0;
    defparam \debounceconsolereset.out_LC_22_10_5 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.out_LC_22_10_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \debounceconsolereset.out_LC_22_10_5  (
            .in0(N__2982),
            .in1(N__2961),
            .in2(N__2940),
            .in3(N__5524),
            .lcout(debouncedconsolereset),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_2_LC_22_11_0.C_ON=1'b0;
    defparam delayConstant_2_LC_22_11_0.SEQ_MODE=4'b1000;
    defparam delayConstant_2_LC_22_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_2_LC_22_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3266),
            .lcout(delayConstantZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5304),
            .ce(),
            .sr(N__4443));
    defparam delayConstant_fast_6_LC_22_11_1.C_ON=1'b0;
    defparam delayConstant_fast_6_LC_22_11_1.SEQ_MODE=4'b1000;
    defparam delayConstant_fast_6_LC_22_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_fast_6_LC_22_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3303),
            .lcout(delayConstant_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5304),
            .ce(),
            .sr(N__4443));
    defparam delayConstant_fast_4_LC_22_11_2.C_ON=1'b0;
    defparam delayConstant_fast_4_LC_22_11_2.SEQ_MODE=4'b1000;
    defparam delayConstant_fast_4_LC_22_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_fast_4_LC_22_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3291),
            .lcout(delayConstant_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5304),
            .ce(),
            .sr(N__4443));
    defparam \arses.counter_0_LC_22_11_3 .C_ON=1'b0;
    defparam \arses.counter_0_LC_22_11_3 .SEQ_MODE=4'b1001;
    defparam \arses.counter_0_LC_22_11_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \arses.counter_0_LC_22_11_3  (
            .in0(_gnd_net_),
            .in1(N__4163),
            .in2(_gnd_net_),
            .in3(N__4556),
            .lcout(\arses.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5304),
            .ce(),
            .sr(N__4443));
    defparam delayConstant_fast_5_LC_22_11_4.C_ON=1'b0;
    defparam delayConstant_fast_5_LC_22_11_4.SEQ_MODE=4'b1001;
    defparam delayConstant_fast_5_LC_22_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 delayConstant_fast_5_LC_22_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3279),
            .lcout(delayConstant_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5304),
            .ce(),
            .sr(N__4443));
    defparam delayConstant_fast_2_LC_22_11_5.C_ON=1'b0;
    defparam delayConstant_fast_2_LC_22_11_5.SEQ_MODE=4'b1000;
    defparam delayConstant_fast_2_LC_22_11_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 delayConstant_fast_2_LC_22_11_5 (
            .in0(N__3267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delayConstant_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5304),
            .ce(),
            .sr(N__4443));
    defparam \dig1.leds_cnst_3_1__m23_bm_LC_22_12_0 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m23_bm_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m23_bm_LC_22_12_0 .LUT_INIT=16'b0100000001110110;
    LogicCell40 \dig1.leds_cnst_3_1__m23_bm_LC_22_12_0  (
            .in0(N__4960),
            .in1(N__3901),
            .in2(N__3466),
            .in3(N__3750),
            .lcout(\dig1.m23_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m8_bm_LC_22_12_6 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m8_bm_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m8_bm_LC_22_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \dig1.leds_cnst_3_1__m8_bm_LC_22_12_6  (
            .in0(N__4959),
            .in1(N__3900),
            .in2(N__3465),
            .in3(N__3751),
            .lcout(\dig1.m8_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m8_am_LC_22_13_0 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m8_am_LC_22_13_0 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m8_am_LC_22_13_0 .LUT_INIT=16'b1101000001111010;
    LogicCell40 \dig1.leds_cnst_3_1__m8_am_LC_22_13_0  (
            .in0(N__4982),
            .in1(N__3906),
            .in2(N__3468),
            .in3(N__3754),
            .lcout(),
            .ltout(\dig1.m8_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m8_ns_LC_22_13_1 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m8_ns_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m8_ns_LC_22_13_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \dig1.leds_cnst_3_1__m8_ns_LC_22_13_1  (
            .in0(N__3373),
            .in1(_gnd_net_),
            .in2(N__3258),
            .in3(N__3255),
            .lcout(),
            .ltout(\dig1.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m13_LC_22_13_2 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m13_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m13_LC_22_13_2 .LUT_INIT=16'b1000110110101111;
    LogicCell40 \dig1.leds_cnst_3_1__m13_LC_22_13_2  (
            .in0(N__4800),
            .in1(N__3519),
            .in2(N__3249),
            .in3(N__3374),
            .lcout(\dig1.leds_cnst_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m11_LC_22_13_3 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m11_LC_22_13_3 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m11_LC_22_13_3 .LUT_INIT=16'b0101011010100101;
    LogicCell40 \dig1.leds_cnst_3_1__m11_LC_22_13_3  (
            .in0(N__3752),
            .in1(N__4980),
            .in2(N__3934),
            .in3(N__3440),
            .lcout(\dig1.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m29_bm_LC_22_13_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m29_bm_LC_22_13_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m29_bm_LC_22_13_4 .LUT_INIT=16'b0100111010110011;
    LogicCell40 \dig1.leds_cnst_3_1__m29_bm_LC_22_13_4  (
            .in0(N__4981),
            .in1(N__3905),
            .in2(N__3467),
            .in3(N__3753),
            .lcout(),
            .ltout(\dig1.m29_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m30_ns_1_LC_22_13_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m30_ns_1_LC_22_13_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m30_ns_1_LC_22_13_5 .LUT_INIT=16'b0000101001110111;
    LogicCell40 \dig1.leds_cnst_3_1__m30_ns_1_LC_22_13_5  (
            .in0(N__3372),
            .in1(N__3513),
            .in2(N__3507),
            .in3(N__4799),
            .lcout(\dig1.m30_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m23_am_LC_22_14_0 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m23_am_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m23_am_LC_22_14_0 .LUT_INIT=16'b1111110001111011;
    LogicCell40 \dig1.leds_cnst_3_1__m23_am_LC_22_14_0  (
            .in0(N__4995),
            .in1(N__3915),
            .in2(N__3487),
            .in3(N__3763),
            .lcout(\dig1.m23_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.un1_leds114_LC_22_14_2 .C_ON=1'b0;
    defparam \dig1.un1_leds114_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \dig1.un1_leds114_LC_22_14_2 .LUT_INIT=16'b1101111111110111;
    LogicCell40 \dig1.un1_leds114_LC_22_14_2  (
            .in0(N__4997),
            .in1(N__3379),
            .in2(N__3489),
            .in3(N__4801),
            .lcout(\dig1.un1_leds114_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m29_am_LC_22_14_4 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m29_am_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m29_am_LC_22_14_4 .LUT_INIT=16'b0000010011111111;
    LogicCell40 \dig1.leds_cnst_3_1__m29_am_LC_22_14_4  (
            .in0(N__4996),
            .in1(N__3916),
            .in2(N__3488),
            .in3(N__3764),
            .lcout(),
            .ltout(\dig1.m29_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m30_ns_LC_22_14_5 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m30_ns_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m30_ns_LC_22_14_5 .LUT_INIT=16'b0100010011111010;
    LogicCell40 \dig1.leds_cnst_3_1__m30_ns_LC_22_14_5  (
            .in0(N__3378),
            .in1(N__3504),
            .in2(N__3498),
            .in3(N__3495),
            .lcout(\dig1.leds_cnst_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_cnst_3_1__m37_LC_22_14_6 .C_ON=1'b0;
    defparam \dig1.leds_cnst_3_1__m37_LC_22_14_6 .SEQ_MODE=4'b0000;
    defparam \dig1.leds_cnst_3_1__m37_LC_22_14_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \dig1.leds_cnst_3_1__m37_LC_22_14_6  (
            .in0(N__3483),
            .in1(N__3917),
            .in2(N__3794),
            .in3(N__3380),
            .lcout(\dig1.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_1_LC_22_15_2 .C_ON=1'b0;
    defparam \dig1.leds_1_i_1_LC_22_15_2 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_1_LC_22_15_2 .LUT_INIT=16'b0101000001010011;
    LogicCell40 \dig1.leds_1_i_1_LC_22_15_2  (
            .in0(N__3333),
            .in1(N__3804),
            .in2(N__4065),
            .in3(N__3947),
            .lcout(leds_1_i_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5309),
            .ce(N__3614),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_3_LC_22_15_3 .C_ON=1'b0;
    defparam \dig1.leds_1_i_3_LC_22_15_3 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_3_LC_22_15_3 .LUT_INIT=16'b1010001100000000;
    LogicCell40 \dig1.leds_1_i_3_LC_22_15_3  (
            .in0(N__4098),
            .in1(N__4092),
            .in2(N__4812),
            .in3(N__4064),
            .lcout(leds_1_i_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5309),
            .ce(N__3614),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_2_LC_22_15_7 .C_ON=1'b0;
    defparam \dig1.leds_1_i_2_LC_22_15_7 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_2_LC_22_15_7 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \dig1.leds_1_i_2_LC_22_15_7  (
            .in0(N__3803),
            .in1(N__4060),
            .in2(_gnd_net_),
            .in3(N__4050),
            .lcout(leds_1_i_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5309),
            .ce(N__3614),
            .sr(_gnd_net_));
    defparam lcolreg_0_LC_22_16_1.C_ON=1'b0;
    defparam lcolreg_0_LC_22_16_1.SEQ_MODE=4'b1000;
    defparam lcolreg_0_LC_22_16_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 lcolreg_0_LC_22_16_1 (
            .in0(_gnd_net_),
            .in1(N__3805),
            .in2(_gnd_net_),
            .in3(N__3946),
            .lcout(lcol1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5310),
            .ce(N__3613),
            .sr(_gnd_net_));
    defparam lcolreg_1_LC_22_17_1.C_ON=1'b0;
    defparam lcolreg_1_LC_22_17_1.SEQ_MODE=4'b1000;
    defparam lcolreg_1_LC_22_17_1.LUT_INIT=16'b1100110011111111;
    LogicCell40 lcolreg_1_LC_22_17_1 (
            .in0(_gnd_net_),
            .in1(N__3948),
            .in2(_gnd_net_),
            .in3(N__3811),
            .lcout(lcol2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5311),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam lcolreg_2_LC_22_17_7.C_ON=1'b0;
    defparam lcolreg_2_LC_22_17_7.SEQ_MODE=4'b1000;
    defparam lcolreg_2_LC_22_17_7.LUT_INIT=16'b1111111100110011;
    LogicCell40 lcolreg_2_LC_22_17_7 (
            .in0(_gnd_net_),
            .in1(N__3949),
            .in2(_gnd_net_),
            .in3(N__3812),
            .lcout(lcol3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5311),
            .ce(N__3627),
            .sr(_gnd_net_));
    defparam lcolreg_3_LC_22_18_5.C_ON=1'b0;
    defparam lcolreg_3_LC_22_18_5.SEQ_MODE=4'b1000;
    defparam lcolreg_3_LC_22_18_5.LUT_INIT=16'b0011001111111111;
    LogicCell40 lcolreg_3_LC_22_18_5 (
            .in0(_gnd_net_),
            .in1(N__3954),
            .in2(_gnd_net_),
            .in3(N__3810),
            .lcout(lcol4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5312),
            .ce(N__3628),
            .sr(_gnd_net_));
    defparam \arse.doingseven_LC_23_7_7 .C_ON=1'b0;
    defparam \arse.doingseven_LC_23_7_7 .SEQ_MODE=4'b1000;
    defparam \arse.doingseven_LC_23_7_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \arse.doingseven_LC_23_7_7  (
            .in0(N__5725),
            .in1(N__4709),
            .in2(_gnd_net_),
            .in3(N__4359),
            .lcout(\arse.doingsevenZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.doingsevenC_net ),
            .ce(),
            .sr(N__5123));
    defparam \arse.cpuresetoutreg_RNO_6_LC_23_8_1 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_6_LC_23_8_1 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_6_LC_23_8_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \arse.cpuresetoutreg_RNO_6_LC_23_8_1  (
            .in0(N__3543),
            .in1(N__3531),
            .in2(N__4674),
            .in3(N__4644),
            .lcout(),
            .ltout(\arse.g0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_3_LC_23_8_2 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_3_LC_23_8_2 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_3_LC_23_8_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \arse.cpuresetoutreg_RNO_3_LC_23_8_2  (
            .in0(_gnd_net_),
            .in1(N__4716),
            .in2(N__4215),
            .in3(N__4830),
            .lcout(),
            .ltout(\arse.g0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_0_LC_23_8_3 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_0_LC_23_8_3 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_0_LC_23_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \arse.cpuresetoutreg_RNO_0_LC_23_8_3  (
            .in0(N__5730),
            .in1(N__4905),
            .in2(N__4212),
            .in3(N__4350),
            .lcout(),
            .ltout(\arse.cpuresetoutreg_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_LC_23_8_4 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_LC_23_8_4 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetoutreg_LC_23_8_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \arse.cpuresetoutreg_LC_23_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4209),
            .in3(N__4196),
            .lcout(\arse.cpuresetoutregZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuresetoutregC_net ),
            .ce(),
            .sr(N__5124));
    defparam \arses.counter_RNIA58_5_LC_23_9_3 .C_ON=1'b0;
    defparam \arses.counter_RNIA58_5_LC_23_9_3 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIA58_5_LC_23_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \arses.counter_RNIA58_5_LC_23_9_3  (
            .in0(N__4283),
            .in1(N__4298),
            .in2(N__4269),
            .in3(N__4313),
            .lcout(),
            .ltout(\arses.un1_counterlto8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOKH_1_LC_23_9_4 .C_ON=1'b0;
    defparam \arses.counter_RNIOKH_1_LC_23_9_4 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOKH_1_LC_23_9_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \arses.counter_RNIOKH_1_LC_23_9_4  (
            .in0(N__4328),
            .in1(N__4133),
            .in2(N__4182),
            .in3(N__4179),
            .lcout(),
            .ltout(\arses.un1_counterlt11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI04C4_9_LC_23_9_5 .C_ON=1'b0;
    defparam \arses.counter_RNI04C4_9_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI04C4_9_LC_23_9_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \arses.counter_RNI04C4_9_LC_23_9_5  (
            .in0(N__4611),
            .in1(N__4233),
            .in2(N__4173),
            .in3(N__4251),
            .lcout(),
            .ltout(\arses.un1_counterlt13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOS0A_14_LC_23_9_6 .C_ON=1'b0;
    defparam \arses.counter_RNIOS0A_14_LC_23_9_6 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOS0A_14_LC_23_9_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \arses.counter_RNIOS0A_14_LC_23_9_6  (
            .in0(N__4593),
            .in1(N__4464),
            .in2(N__4170),
            .in3(N__4575),
            .lcout(\arses.counter8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.un2_counter_cry_1_c_LC_23_10_0 .C_ON=1'b1;
    defparam \arses.un2_counter_cry_1_c_LC_23_10_0 .SEQ_MODE=4'b0000;
    defparam \arses.un2_counter_cry_1_c_LC_23_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \arses.un2_counter_cry_1_c_LC_23_10_0  (
            .in0(_gnd_net_),
            .in1(N__4162),
            .in2(N__4140),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_23_10_0_),
            .carryout(\arses.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_2_LC_23_10_1 .C_ON=1'b1;
    defparam \arses.counter_2_LC_23_10_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_2_LC_23_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_2_LC_23_10_1  (
            .in0(N__4551),
            .in1(N__4113),
            .in2(_gnd_net_),
            .in3(N__4101),
            .lcout(\arses.counterZ0Z_2 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_1 ),
            .carryout(\arses.un2_counter_cry_2 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_3_LC_23_10_2 .C_ON=1'b1;
    defparam \arses.counter_3_LC_23_10_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_3_LC_23_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_3_LC_23_10_2  (
            .in0(N__4533),
            .in1(N__4344),
            .in2(_gnd_net_),
            .in3(N__4332),
            .lcout(\arses.counterZ0Z_3 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_2 ),
            .carryout(\arses.un2_counter_cry_3 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_4_LC_23_10_3 .C_ON=1'b1;
    defparam \arses.counter_4_LC_23_10_3 .SEQ_MODE=4'b1001;
    defparam \arses.counter_4_LC_23_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_4_LC_23_10_3  (
            .in0(N__4552),
            .in1(N__4329),
            .in2(_gnd_net_),
            .in3(N__4317),
            .lcout(\arses.counterZ0Z_4 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_3 ),
            .carryout(\arses.un2_counter_cry_4 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_5_LC_23_10_4 .C_ON=1'b1;
    defparam \arses.counter_5_LC_23_10_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_5_LC_23_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_5_LC_23_10_4  (
            .in0(N__4534),
            .in1(N__4314),
            .in2(_gnd_net_),
            .in3(N__4302),
            .lcout(\arses.counterZ0Z_5 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_4 ),
            .carryout(\arses.un2_counter_cry_5 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_6_LC_23_10_5 .C_ON=1'b1;
    defparam \arses.counter_6_LC_23_10_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_6_LC_23_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_6_LC_23_10_5  (
            .in0(N__4553),
            .in1(N__4299),
            .in2(_gnd_net_),
            .in3(N__4287),
            .lcout(\arses.counterZ0Z_6 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_5 ),
            .carryout(\arses.un2_counter_cry_6 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_7_LC_23_10_6 .C_ON=1'b1;
    defparam \arses.counter_7_LC_23_10_6 .SEQ_MODE=4'b1000;
    defparam \arses.counter_7_LC_23_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_7_LC_23_10_6  (
            .in0(N__4535),
            .in1(N__4284),
            .in2(_gnd_net_),
            .in3(N__4272),
            .lcout(\arses.counterZ0Z_7 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_6 ),
            .carryout(\arses.un2_counter_cry_7 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_8_LC_23_10_7 .C_ON=1'b1;
    defparam \arses.counter_8_LC_23_10_7 .SEQ_MODE=4'b1000;
    defparam \arses.counter_8_LC_23_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_8_LC_23_10_7  (
            .in0(N__4554),
            .in1(N__4268),
            .in2(_gnd_net_),
            .in3(N__4254),
            .lcout(\arses.counterZ0Z_8 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_7 ),
            .carryout(\arses.un2_counter_cry_8 ),
            .clk(N__5305),
            .ce(),
            .sr(N__4446));
    defparam \arses.counter_9_LC_23_11_0 .C_ON=1'b1;
    defparam \arses.counter_9_LC_23_11_0 .SEQ_MODE=4'b1000;
    defparam \arses.counter_9_LC_23_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_9_LC_23_11_0  (
            .in0(N__4547),
            .in1(N__4250),
            .in2(_gnd_net_),
            .in3(N__4236),
            .lcout(\arses.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_23_11_0_),
            .carryout(\arses.un2_counter_cry_9 ),
            .clk(N__5307),
            .ce(),
            .sr(N__4445));
    defparam \arses.counter_10_LC_23_11_1 .C_ON=1'b1;
    defparam \arses.counter_10_LC_23_11_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_10_LC_23_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_10_LC_23_11_1  (
            .in0(N__4548),
            .in1(N__4232),
            .in2(_gnd_net_),
            .in3(N__4218),
            .lcout(\arses.counterZ0Z_10 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_9 ),
            .carryout(\arses.un2_counter_cry_10 ),
            .clk(N__5307),
            .ce(),
            .sr(N__4445));
    defparam \arses.counter_11_LC_23_11_2 .C_ON=1'b1;
    defparam \arses.counter_11_LC_23_11_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_11_LC_23_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_11_LC_23_11_2  (
            .in0(N__4545),
            .in1(N__4610),
            .in2(_gnd_net_),
            .in3(N__4596),
            .lcout(\arses.counterZ0Z_11 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_10 ),
            .carryout(\arses.un2_counter_cry_11 ),
            .clk(N__5307),
            .ce(),
            .sr(N__4445));
    defparam \arses.counter_12_LC_23_11_3 .C_ON=1'b1;
    defparam \arses.counter_12_LC_23_11_3 .SEQ_MODE=4'b1000;
    defparam \arses.counter_12_LC_23_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_12_LC_23_11_3  (
            .in0(N__4549),
            .in1(N__4592),
            .in2(_gnd_net_),
            .in3(N__4578),
            .lcout(\arses.counterZ0Z_12 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_11 ),
            .carryout(\arses.un2_counter_cry_12 ),
            .clk(N__5307),
            .ce(),
            .sr(N__4445));
    defparam \arses.counter_13_LC_23_11_4 .C_ON=1'b1;
    defparam \arses.counter_13_LC_23_11_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_13_LC_23_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_13_LC_23_11_4  (
            .in0(N__4546),
            .in1(N__4574),
            .in2(_gnd_net_),
            .in3(N__4560),
            .lcout(\arses.counterZ0Z_13 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_12 ),
            .carryout(\arses.un2_counter_cry_13 ),
            .clk(N__5307),
            .ce(),
            .sr(N__4445));
    defparam \arses.counter_14_LC_23_11_5 .C_ON=1'b0;
    defparam \arses.counter_14_LC_23_11_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_14_LC_23_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_14_LC_23_11_5  (
            .in0(N__4550),
            .in1(N__4460),
            .in2(_gnd_net_),
            .in3(N__4467),
            .lcout(\arses.counterZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5307),
            .ce(),
            .sr(N__4445));
    defparam CONSTANT_ONE_LUT4_LC_23_31_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_23_31_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_23_31_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_23_31_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.doingseven_RNO_0_LC_24_7_1 .C_ON=1'b0;
    defparam \arse.doingseven_RNO_0_LC_24_7_1 .SEQ_MODE=4'b0000;
    defparam \arse.doingseven_RNO_0_LC_24_7_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \arse.doingseven_RNO_0_LC_24_7_1  (
            .in0(N__4686),
            .in1(N__4647),
            .in2(N__4695),
            .in3(N__4739),
            .lcout(\arse.doingseven3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_RNIB4QP_0_LC_24_7_3 .C_ON=1'b0;
    defparam \arse.cpuresetcount_RNIB4QP_0_LC_24_7_3 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetcount_RNIB4QP_0_LC_24_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.cpuresetcount_RNIB4QP_0_LC_24_7_3  (
            .in0(_gnd_net_),
            .in1(N__4668),
            .in2(_gnd_net_),
            .in3(N__5022),
            .lcout(\arse.doingseven3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_4_LC_24_7_4 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_4_LC_24_7_4 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_4_LC_24_7_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \arse.cpuresetoutreg_RNO_4_LC_24_7_4  (
            .in0(N__4669),
            .in1(N__4759),
            .in2(N__5025),
            .in3(N__4849),
            .lcout(),
            .ltout(\arse.g0_i_a3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_1_LC_24_7_5 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_1_LC_24_7_5 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_1_LC_24_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \arse.cpuresetoutreg_RNO_1_LC_24_7_5  (
            .in0(N__4929),
            .in1(N__4870),
            .in2(N__4353),
            .in3(N__4737),
            .lcout(\arse.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_RNIATKJ1_7_LC_24_7_6 .C_ON=1'b0;
    defparam \arse.cpuresetcount_RNIATKJ1_7_LC_24_7_6 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetcount_RNIATKJ1_7_LC_24_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \arse.cpuresetcount_RNIATKJ1_7_LC_24_7_6  (
            .in0(N__4869),
            .in1(N__4758),
            .in2(N__4932),
            .in3(N__4850),
            .lcout(\arse.doingseven3_6 ),
            .ltout(\arse.doingseven3_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuclkreset_RNO_0_LC_24_7_7 .C_ON=1'b0;
    defparam \arse.cpuclkreset_RNO_0_LC_24_7_7 .SEQ_MODE=4'b0000;
    defparam \arse.cpuclkreset_RNO_0_LC_24_7_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \arse.cpuclkreset_RNO_0_LC_24_7_7  (
            .in0(N__4685),
            .in1(N__4646),
            .in2(N__4677),
            .in3(N__4738),
            .lcout(\arse.doingseven4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_0_LC_24_8_0 .C_ON=1'b1;
    defparam \arse.cpuresetcount_0_LC_24_8_0 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_0_LC_24_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_0_LC_24_8_0  (
            .in0(_gnd_net_),
            .in1(N__4670),
            .in2(N__5729),
            .in3(N__5724),
            .lcout(\arse.cpuresetcountZ0Z_0 ),
            .ltout(),
            .carryin(bfn_24_8_0_),
            .carryout(\arse.un1_cpuresetcount_1_cry_0 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_1_LC_24_8_1 .C_ON=1'b1;
    defparam \arse.cpuresetcount_1_LC_24_8_1 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_1_LC_24_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_1_LC_24_8_1  (
            .in0(_gnd_net_),
            .in1(N__5024),
            .in2(_gnd_net_),
            .in3(N__4650),
            .lcout(\arse.cpuresetcountZ0Z_1 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_0 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_1 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_2_LC_24_8_2 .C_ON=1'b1;
    defparam \arse.cpuresetcount_2_LC_24_8_2 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_2_LC_24_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_2_LC_24_8_2  (
            .in0(_gnd_net_),
            .in1(N__4645),
            .in2(_gnd_net_),
            .in3(N__4626),
            .lcout(\arse.cpuresetcountZ0Z_2 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_1 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_2 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_3_LC_24_8_3 .C_ON=1'b1;
    defparam \arse.cpuresetcount_3_LC_24_8_3 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_3_LC_24_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_3_LC_24_8_3  (
            .in0(_gnd_net_),
            .in1(N__4740),
            .in2(_gnd_net_),
            .in3(N__4623),
            .lcout(\arse.cpuresetcountZ0Z_3 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_2 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_3 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_4_LC_24_8_4 .C_ON=1'b1;
    defparam \arse.cpuresetcount_4_LC_24_8_4 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_4_LC_24_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_4_LC_24_8_4  (
            .in0(_gnd_net_),
            .in1(N__4763),
            .in2(_gnd_net_),
            .in3(N__4620),
            .lcout(\arse.cpuresetcountZ0Z_4 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_3 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_4 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_5_LC_24_8_5 .C_ON=1'b1;
    defparam \arse.cpuresetcount_5_LC_24_8_5 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_5_LC_24_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_5_LC_24_8_5  (
            .in0(_gnd_net_),
            .in1(N__4851),
            .in2(_gnd_net_),
            .in3(N__4617),
            .lcout(\arse.cpuresetcountZ0Z_5 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_4 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_5 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_6_LC_24_8_6 .C_ON=1'b1;
    defparam \arse.cpuresetcount_6_LC_24_8_6 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_6_LC_24_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_6_LC_24_8_6  (
            .in0(_gnd_net_),
            .in1(N__4874),
            .in2(_gnd_net_),
            .in3(N__4614),
            .lcout(\arse.cpuresetcountZ0Z_6 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_5 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_6 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetcount_7_LC_24_8_7 .C_ON=1'b0;
    defparam \arse.cpuresetcount_7_LC_24_8_7 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_7_LC_24_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \arse.cpuresetcount_7_LC_24_8_7  (
            .in0(_gnd_net_),
            .in1(N__4931),
            .in2(_gnd_net_),
            .in3(N__5079),
            .lcout(\arse.cpuresetcountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5115));
    defparam \arse.cpuresetoutreg_RNO_2_LC_24_9_4 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_2_LC_24_9_4 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_2_LC_24_9_4 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \arse.cpuresetoutreg_RNO_2_LC_24_9_4  (
            .in0(N__5075),
            .in1(N__5023),
            .in2(N__5001),
            .in3(N__4930),
            .lcout(\arse.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_7_LC_24_9_6 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_7_LC_24_9_6 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_7_LC_24_9_6 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \arse.cpuresetoutreg_RNO_7_LC_24_9_6  (
            .in0(N__4899),
            .in1(N__4887),
            .in2(N__4875),
            .in3(N__4848),
            .lcout(\arse.g0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_5_LC_24_9_7 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_5_LC_24_9_7 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_5_LC_24_9_7 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \arse.cpuresetoutreg_RNO_5_LC_24_9_7  (
            .in0(N__4824),
            .in1(N__4811),
            .in2(N__4764),
            .in3(N__4736),
            .lcout(\arse.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.seven_LC_26_7_6 .C_ON=1'b0;
    defparam \arse.divseven.seven_LC_26_7_6 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.seven_LC_26_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.divseven.seven_LC_26_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4710),
            .lcout(\arse.divseven.sevenZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5391),
            .ce(N__5352),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_2_LC_26_8_0 .C_ON=1'b0;
    defparam \arse.divseven.counter_2_LC_26_8_0 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_2_LC_26_8_0 .LUT_INIT=16'b1001111110100000;
    LogicCell40 \arse.divseven.counter_2_LC_26_8_0  (
            .in0(N__5437),
            .in1(N__5161),
            .in2(N__5196),
            .in3(N__5492),
            .lcout(\arse.divseven.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5390),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_0_LC_26_8_2 .C_ON=1'b0;
    defparam \arse.divseven.counter_0_LC_26_8_2 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_0_LC_26_8_2 .LUT_INIT=16'b1001010101010101;
    LogicCell40 \arse.divseven.counter_0_LC_26_8_2  (
            .in0(N__5436),
            .in1(N__5157),
            .in2(N__5195),
            .in3(N__5491),
            .lcout(\arse.divseven.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5390),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_1_LC_26_8_3 .C_ON=1'b0;
    defparam \arse.divseven.counter_1_LC_26_8_3 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_1_LC_26_8_3 .LUT_INIT=16'b1011001101001100;
    LogicCell40 \arse.divseven.counter_1_LC_26_8_3  (
            .in0(N__5490),
            .in1(N__5187),
            .in2(N__5163),
            .in3(N__5438),
            .lcout(\arse.divseven.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5390),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.seven_RNO_LC_26_8_5 .C_ON=1'b0;
    defparam \arse.divseven.seven_RNO_LC_26_8_5 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.seven_RNO_LC_26_8_5 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \arse.divseven.seven_RNO_LC_26_8_5  (
            .in0(N__5489),
            .in1(N__5186),
            .in2(N__5162),
            .in3(N__5435),
            .lcout(\arse.divseven.N_41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.out_e_0_LC_26_10_5 .C_ON=1'b0;
    defparam \debounceup.out_e_0_LC_26_10_5 .SEQ_MODE=4'b1000;
    defparam \debounceup.out_e_0_LC_26_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceup.out_e_0_LC_26_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5340),
            .lcout(debouncedup),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5308),
            .ce(N__5241),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_RNO_0_0_LC_27_8_2 .C_ON=1'b0;
    defparam \arse.divseven.dout_RNO_0_0_LC_27_8_2 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.dout_RNO_0_0_LC_27_8_2 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \arse.divseven.dout_RNO_0_0_LC_27_8_2  (
            .in0(N__5434),
            .in1(N__5207),
            .in2(N__5194),
            .in3(N__5487),
            .lcout(),
            .ltout(\arse.divseven.dout_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_0_LC_27_8_3 .C_ON=1'b0;
    defparam \arse.divseven.dout_0_LC_27_8_3 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_0_LC_27_8_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \arse.divseven.dout_0_LC_27_8_3  (
            .in0(N__5488),
            .in1(_gnd_net_),
            .in2(N__5220),
            .in3(N__5152),
            .lcout(\arse.divseven.doutZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.divseven.dout_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_RNO_0_1_LC_27_8_7 .C_ON=1'b0;
    defparam \arse.divseven.dout_RNO_0_1_LC_27_8_7 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.dout_RNO_0_1_LC_27_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.divseven.dout_RNO_0_1_LC_27_8_7  (
            .in0(_gnd_net_),
            .in1(N__5185),
            .in2(_gnd_net_),
            .in3(N__5153),
            .lcout(\arse.divseven.un1_dout_2_sqmuxa_0_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_1 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \debounceconsolereset.out_RNI1B6C_LC_29_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5548),
            .lcout(debouncedconsolereset_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuclkreset_LC_30_7_6 .C_ON=1'b0;
    defparam \arse.cpuclkreset_LC_30_7_6 .SEQ_MODE=4'b1000;
    defparam \arse.cpuclkreset_LC_30_7_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \arse.cpuclkreset_LC_30_7_6  (
            .in0(N__5698),
            .in1(N__5614),
            .in2(_gnd_net_),
            .in3(N__5133),
            .lcout(\arse.cpuclkresetZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuclkresetC_net ),
            .ce(),
            .sr(N__5122));
    defparam \arse.diveight.counter_2_LC_31_6_1 .C_ON=1'b0;
    defparam \arse.diveight.counter_2_LC_31_6_1 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_2_LC_31_6_1 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \arse.diveight.counter_2_LC_31_6_1  (
            .in0(N__5671),
            .in1(N__5607),
            .in2(N__5648),
            .in3(N__5579),
            .lcout(\arse.diveight.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_0_LC_31_6_5 .C_ON=1'b0;
    defparam \arse.diveight.counter_0_LC_31_6_5 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_0_LC_31_6_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \arse.diveight.counter_0_LC_31_6_5  (
            .in0(_gnd_net_),
            .in1(N__5667),
            .in2(_gnd_net_),
            .in3(N__5605),
            .lcout(\arse.diveight.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_1_LC_31_6_6 .C_ON=1'b0;
    defparam \arse.diveight.counter_1_LC_31_6_6 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_1_LC_31_6_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \arse.diveight.counter_1_LC_31_6_6  (
            .in0(N__5606),
            .in1(_gnd_net_),
            .in2(N__5673),
            .in3(N__5641),
            .lcout(\arse.diveight.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5396),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.apusynclatched_LC_32_4_3 .C_ON=1'b0;
    defparam \arse.apusynclatched_LC_32_4_3 .SEQ_MODE=4'b1000;
    defparam \arse.apusynclatched_LC_32_4_3 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \arse.apusynclatched_LC_32_4_3  (
            .in0(N__5742),
            .in1(N__5684),
            .in2(_gnd_net_),
            .in3(N__5556),
            .lcout(\arse.apusynclatchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.apusynclatchedC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_1_LC_32_5_0 .C_ON=1'b0;
    defparam \arse.diveight.dout_1_LC_32_5_0 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_1_LC_32_5_0 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \arse.diveight.dout_1_LC_32_5_0  (
            .in0(N__5672),
            .in1(N__5621),
            .in2(N__5649),
            .in3(N__5580),
            .lcout(\arse.diveight.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5398),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_0_LC_32_6_5 .C_ON=1'b0;
    defparam \arse.diveight.dout_0_LC_32_6_5 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_0_LC_32_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.diveight.dout_0_LC_32_6_5  (
            .in0(_gnd_net_),
            .in1(N__5622),
            .in2(_gnd_net_),
            .in3(N__5578),
            .lcout(\arse.diveight.doutZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.diveight.dout_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.apuresetoutreg_LC_32_6_6 .C_ON=1'b0;
    defparam \arse.apuresetoutreg_LC_32_6_6 .SEQ_MODE=4'b1000;
    defparam \arse.apuresetoutreg_LC_32_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.apuresetoutreg_LC_32_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5555),
            .lcout(\arse.apuresetoutregZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.diveight.dout_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_1_LC_32_9_4 .C_ON=1'b0;
    defparam \arse.divseven.dout_1_LC_32_9_4 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_1_LC_32_9_4 .LUT_INIT=16'b1011110011001100;
    LogicCell40 \arse.divseven.dout_1_LC_32_9_4  (
            .in0(N__5412),
            .in1(N__5502),
            .in2(N__5463),
            .in3(N__5445),
            .lcout(\arse.divseven.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5394),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
