-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 11 2024 23:52:07

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    masterreset : in std_logic;
    led4 : out std_logic;
    lcol3 : out std_logic;
    led5 : out std_logic;
    lcol2 : out std_logic;
    led6 : out std_logic;
    led2 : out std_logic;
    lcol1 : out std_logic;
    deldn : in std_logic;
    cpuclk : out std_logic;
    apureset : out std_logic;
    led7 : out std_logic;
    led3 : out std_logic;
    lcol4 : out std_logic;
    delup : in std_logic;
    cpureset : out std_logic;
    apusync : in std_logic;
    PACKAGEPIN : in std_logic;
    led8 : out std_logic;
    led1 : out std_logic;
    consolereset : in std_logic;
    apuclk : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \arse.un1_io_0_1_g\ : std_logic;
signal \top_pll_nrtthrth.PLLOUTCORE\ : std_logic;
signal \GNDG0\ : std_logic;
signal \arse.divseven.io_0_D_IN_0\ : std_logic;
signal \VCCG0\ : std_logic;
signal masterreset_c_i : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \debouncedn.un3_counter_cry_1\ : std_logic;
signal \debouncedn.un3_counter_cry_2\ : std_logic;
signal \debouncedn.un3_counter_cry_3\ : std_logic;
signal \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\ : std_logic;
signal \debouncedn.counter18_0_2_cascade_\ : std_logic;
signal \debouncedn.counterZ0Z_1\ : std_logic;
signal \debouncedn.counterZ0Z_4\ : std_logic;
signal \debouncedn.counter_RNIBTPA2Z0Z_4_cascade_\ : std_logic;
signal \debouncedn.counterZ0Z_0\ : std_logic;
signal \debounceconsolereset.counter18_0_2_cascade_\ : std_logic;
signal \debouncedn.un3_counter_cry_2_THRU_CO\ : std_logic;
signal \debouncedn.counterZ0Z_3\ : std_logic;
signal \debouncedn.un3_counter_cry_1_THRU_CO\ : std_logic;
signal \debouncedn.counter_RNIBTPA2Z0Z_4\ : std_logic;
signal \debouncedn.counterZ0Z_2\ : std_logic;
signal consolereset_c : std_logic;
signal \debounceconsolereset.out_cnv_2\ : std_logic;
signal lcol3_c : std_logic;
signal lcol4_c : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \debounceup.un3_counter_cry_1\ : std_logic;
signal \debounceup.un3_counter_cry_2\ : std_logic;
signal \debounceup.un3_counter_cry_3\ : std_logic;
signal \debounceup.un3_counter_cry_2_THRU_CO\ : std_logic;
signal \debounceup.un3_counter_cry_1_THRU_CO\ : std_logic;
signal \debounceconsolereset.counterZ0Z_1\ : std_logic;
signal \debounceconsolereset.counterZ0Z_0\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_1\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_2\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_3\ : std_logic;
signal \debounceconsolereset.counterZ0Z_4\ : std_logic;
signal \clock_out_RNIR6ER_0_cascade_\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_2_THRU_CO\ : std_logic;
signal \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_\ : std_logic;
signal \debounceconsolereset.counterZ0Z_3\ : std_logic;
signal \debounceconsolereset.counter_RNINST81Z0Z_4\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_1_THRU_CO\ : std_logic;
signal \debounceconsolereset.counterZ0Z_2\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \arses.un2_counter_cry_1\ : std_logic;
signal \arses.un2_counter_cry_2\ : std_logic;
signal \arses.un2_counter_cry_3\ : std_logic;
signal \arses.un2_counter_cry_4\ : std_logic;
signal \arses.un2_counter_cry_5\ : std_logic;
signal \arses.un2_counter_cry_6\ : std_logic;
signal \arses.un2_counter_cry_7\ : std_logic;
signal \arses.un2_counter_cry_8\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \arses.un2_counter_cry_9\ : std_logic;
signal \arses.un2_counter_cry_10\ : std_logic;
signal \arses.un2_counter_cry_11\ : std_logic;
signal \arses.un2_counter_cry_12\ : std_logic;
signal \arses.un2_counter_cry_13\ : std_logic;
signal leds_1_i_0_3 : std_logic;
signal \debounceup.counter_RNI45V02Z0Z_4_cascade_\ : std_logic;
signal \debounceup.counterZ0Z_3\ : std_logic;
signal \debounceup.counterZ0Z_2\ : std_logic;
signal \debounceup.counterZ0Z_4\ : std_logic;
signal \debounceup.counter18_0_2_cascade_\ : std_logic;
signal \debounceup.counterZ0Z_0\ : std_logic;
signal \debounceup.counter_RNI45V02Z0Z_4\ : std_logic;
signal \debounceup.counterZ0Z_1\ : std_logic;
signal leds_1_i_0_2 : std_logic;
signal \arses.counterZ0Z_7\ : std_logic;
signal \arses.counterZ0Z_6\ : std_logic;
signal \arses.counterZ0Z_8\ : std_logic;
signal \arses.counterZ0Z_5\ : std_logic;
signal \arses.counterZ0Z_4\ : std_logic;
signal \arses.counterZ0Z_1\ : std_logic;
signal \arses.un1_counterlto8_2_cascade_\ : std_logic;
signal \arses.counterZ0Z_11\ : std_logic;
signal \arses.counterZ0Z_10\ : std_logic;
signal \arses.un1_counterlt11_cascade_\ : std_logic;
signal \arses.counterZ0Z_9\ : std_logic;
signal \arses.counterZ0Z_14\ : std_logic;
signal \arses.counterZ0Z_13\ : std_logic;
signal \arses.un1_counterlt13_0_cascade_\ : std_logic;
signal \arses.counterZ0Z_12\ : std_logic;
signal \arses.counter8_cascade_\ : std_logic;
signal \arses.counterZ0Z_3\ : std_logic;
signal \arses.counterZ0Z_2\ : std_logic;
signal \arses.un1_counterlto4_2\ : std_logic;
signal \arses.counterZ0Z_0\ : std_logic;
signal \dig1.N_78\ : std_logic;
signal \dig1.N_72\ : std_logic;
signal \debouncedn.out_cnv_2\ : std_logic;
signal deldn_c : std_logic;
signal \dig1.N_58_cascade_\ : std_logic;
signal \dig1.leds_17_i_ns_1_2\ : std_logic;
signal \dig1.N_61\ : std_logic;
signal \dig1.m68_bm\ : std_logic;
signal \dig1.m68_am\ : std_logic;
signal \arses.counter8\ : std_logic;
signal lcol2_c : std_logic;
signal masterreset_c : std_logic;
signal \delayConstant16_i_cascade_\ : std_logic;
signal \oldupZ0\ : std_logic;
signal debounceddn : std_logic;
signal \olddnZ0\ : std_logic;
signal \dig1.m77_am\ : std_logic;
signal \debounceup.out_cnv_2\ : std_logic;
signal delup_c : std_logic;
signal debouncedup : std_logic;
signal \dig1.m77_bm\ : std_logic;
signal leds_1_i_1 : std_logic;
signal lcol1_c : std_logic;
signal \dig1.N_39\ : std_logic;
signal leds_1_i_3 : std_logic;
signal \dig1.N_15_cascade_\ : std_logic;
signal \dig1.N_18\ : std_logic;
signal slowclk : std_logic;
signal \clock_out_RNIR6ER\ : std_logic;
signal \dig1.N_17\ : std_logic;
signal \dig1.m32_bm\ : std_logic;
signal \dig1.m32_am\ : std_logic;
signal leds_1_i_2 : std_logic;
signal \un1_delayConstant_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_21_12_0_\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_1\ : std_logic;
signal \un1_delayConstant_cry_0\ : std_logic;
signal \olddn_RNIM5BHZ0Z1\ : std_logic;
signal \un1_delayConstant_cry_1\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_2\ : std_logic;
signal \un1_delayConstant_cry_2\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_3\ : std_logic;
signal \un1_delayConstant_cry_3\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_0\ : std_logic;
signal \un1_delayConstant_cry_4\ : std_logic;
signal \olddn_RNIM5BH1Z0Z_4\ : std_logic;
signal \un1_delayConstant_cry_5\ : std_logic;
signal \delayConstant16_i\ : std_logic;
signal \olddn_RNIEENHZ0\ : std_logic;
signal \un1_delayConstant_cry_6\ : std_logic;
signal \dig1.m41_bm\ : std_logic;
signal \dig1.m41_am_cascade_\ : std_logic;
signal \dig1.N_44\ : std_logic;
signal \dig1.m10_ns_1_cascade_\ : std_logic;
signal \dig1.N_11_0\ : std_logic;
signal \delayConstantZ0Z_6\ : std_logic;
signal \dig1.N_25\ : std_logic;
signal \dig1.N_22_cascade_\ : std_logic;
signal \dig1.leds_17_i_0_ns_1_2\ : std_logic;
signal \un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2\ : std_logic;
signal \un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92\ : std_logic;
signal masterreset_c_i_g : std_logic;
signal leds_1_i_0_1 : std_logic;
signal \PACKAGEPIN_0_c_g\ : std_logic;
signal \clock_out_RNIR6ER_0\ : std_logic;
signal \dig1.N_52_cascade_\ : std_logic;
signal \dig1.N_54\ : std_logic;
signal \dig1.N_55\ : std_logic;
signal \colZ0Z_0\ : std_logic;
signal \colZ0Z_1\ : std_logic;
signal \delayConstantZ0Z_2\ : std_logic;
signal \dig1.m47_ns_1_cascade_\ : std_logic;
signal col_1_1 : std_logic;
signal \dig1.N_49\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bfn_27_8_0_\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_0\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_1\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_2\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_3\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_4\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_5\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_6\ : std_logic;
signal \INVarse.cpuresetcount_0C_net\ : std_logic;
signal \delayConstantZ0Z_1\ : std_logic;
signal \delayConstantZ0Z_5\ : std_logic;
signal \arse.g0_i_a3_4\ : std_logic;
signal \arse.cpuresetcountZ0Z_5\ : std_logic;
signal \arse.doingseven3_6_cascade_\ : std_logic;
signal \arse.cpuresetcountZ0Z_1\ : std_logic;
signal \arse.doingseven3_1\ : std_logic;
signal \arse.doingseven3_6\ : std_logic;
signal \arse.doingseven3_1_cascade_\ : std_logic;
signal \delayConstant_fastZ0Z_6\ : std_logic;
signal \delayConstant_fastZ0Z_2\ : std_logic;
signal \arse.cpuresetcountZ0Z_6\ : std_logic;
signal \arse.cpuresetcountZ0Z_2\ : std_logic;
signal \delayConstantZ0Z_7\ : std_logic;
signal \delayConstantZ0Z_3\ : std_logic;
signal \arse.cpuresetcountZ0Z_7\ : std_logic;
signal \arse.cpuresetcountZ0Z_3\ : std_logic;
signal \delayConstantZ0Z_4\ : std_logic;
signal \delayConstantZ0Z_0\ : std_logic;
signal \arse.cpuresetcountZ0Z_0\ : std_logic;
signal \arse.cpuresetcountZ0Z_4\ : std_logic;
signal \arse.g0_3\ : std_logic;
signal \arse.g0_2_cascade_\ : std_logic;
signal \arse.g0_4\ : std_logic;
signal \arse.N_6\ : std_logic;
signal \arse.g0_1\ : std_logic;
signal \arse.g0_7_cascade_\ : std_logic;
signal \arse.cpuresetoutreg_1_sqmuxa_cascade_\ : std_logic;
signal \arse.cpuresetoutregZ0\ : std_logic;
signal \INVarse.cpuresetoutregC_net\ : std_logic;
signal \arse.doingseven4\ : std_logic;
signal \INVarse.cpuclkresetC_net\ : std_logic;
signal \arse.doingseven3\ : std_logic;
signal \INVarse.doingsevenC_net\ : std_logic;
signal debouncedconsolereset_i : std_logic;
signal \arse.doingsevenZ0\ : std_logic;
signal \arse.diveight.doutZ1Z_0\ : std_logic;
signal \INVarse.diveight.dout_0C_net\ : std_logic;
signal \arse.divseven.un1_counter_i_0_0\ : std_logic;
signal \arse.divseven.counterZ0Z_0\ : std_logic;
signal \arse.divseven.sevenZ0\ : std_logic;
signal apusync_c : std_logic;
signal \arse.apusynclatchedZ0\ : std_logic;
signal \INVarse.apusynclatchedC_net\ : std_logic;
signal debouncedconsolereset : std_logic;
signal \arse.apuresetoutregZ0\ : std_logic;
signal \INVarse.apuresetoutregC_net\ : std_logic;
signal \arse.diveight.counterZ0Z_0\ : std_logic;
signal \arse.cpuclkresetZ0\ : std_logic;
signal \arse.diveight.counterZ0Z_1\ : std_logic;
signal \arse.diveight.counterZ0Z_2\ : std_logic;
signal \arse.diveight.doutZ0Z_1\ : std_logic;
signal \arse.divseven.N_46_0\ : std_logic;
signal \arse.divseven.counterZ0Z_1\ : std_logic;
signal \arse.divseven.doutZ0Z_1\ : std_logic;
signal \PLLOUTCORE_g\ : std_logic;
signal \arse.divseven.counterZ0Z_2\ : std_logic;
signal \arse.divseven.doutZ0Z_0\ : std_logic;
signal \INVarse.divseven.dout_0C_net\ : std_logic;
signal \arse.divseven.un1_dout_2_sqmuxa_0_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PACKAGEPIN_wire\ : std_logic;
signal masterreset_wire : std_logic;
signal led3_wire : std_logic;
signal apuclk_wire : std_logic;
signal cpureset_wire : std_logic;
signal lcol3_wire : std_logic;
signal deldn_wire : std_logic;
signal led2_wire : std_logic;
signal delup_wire : std_logic;
signal led6_wire : std_logic;
signal led8_wire : std_logic;
signal led4_wire : std_logic;
signal apureset_wire : std_logic;
signal lcol4_wire : std_logic;
signal cpuclk_wire : std_logic;
signal led5_wire : std_logic;
signal consolereset_wire : std_logic;
signal lcol2_wire : std_logic;
signal led1_wire : std_logic;
signal apusync_wire : std_logic;
signal led7_wire : std_logic;
signal lcol1_wire : std_logic;
signal \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \PACKAGEPIN_wire\ <= PACKAGEPIN;
    masterreset_wire <= masterreset;
    led3 <= led3_wire;
    apuclk <= apuclk_wire;
    cpureset <= cpureset_wire;
    lcol3 <= lcol3_wire;
    deldn_wire <= deldn;
    led2 <= led2_wire;
    delup_wire <= delup;
    led6 <= led6_wire;
    led8 <= led8_wire;
    led4 <= led4_wire;
    apureset <= apureset_wire;
    lcol4 <= lcol4_wire;
    cpuclk <= cpuclk_wire;
    led5 <= led5_wire;
    consolereset_wire <= consolereset;
    lcol2 <= lcol2_wire;
    led1 <= led1_wire;
    apusync_wire <= apusync;
    led7 <= led7_wire;
    lcol1 <= lcol1_wire;
    \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_nrtthrth.top_pll_nrtthrth_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "010",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \top_pll_nrtthrth.PLLOUTCORE\,
            REFERENCECLK => \N__2510\,
            RESETB => \N__3602\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PACKAGEPIN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6474\,
            GLOBALBUFFEROUTPUT => \PACKAGEPIN_0_c_g\
        );

    \PACKAGEPIN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6476\,
            DIN => \N__6475\,
            DOUT => \N__6474\,
            PACKAGEPIN => \PACKAGEPIN_wire\
        );

    \PACKAGEPIN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6476\,
            PADOUT => \N__6475\,
            PADIN => \N__6474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \masterreset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6465\,
            DIN => \N__6464\,
            DOUT => \N__6463\,
            PACKAGEPIN => masterreset_wire
        );

    \masterreset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6465\,
            PADOUT => \N__6464\,
            PADIN => \N__6463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => masterreset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6456\,
            DIN => \N__6455\,
            DOUT => \N__6454\,
            PACKAGEPIN => led3_wire
        );

    \led3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6456\,
            PADOUT => \N__6455\,
            PADIN => \N__6454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.divseven.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6447\,
            DIN => \N__6446\,
            DOUT => \N__6445\,
            PACKAGEPIN => apuclk_wire
        );

    \arse.divseven.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6447\,
            PADOUT => \N__6446\,
            PADIN => \N__6445\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__5926\,
            OUTPUTENABLE => \N__4973\,
            DIN0 => \arse.divseven.io_0_D_IN_0\,
            DOUT0 => \N__5834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5909\
        );

    \arse.io_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6438\,
            DIN => \N__6437\,
            DOUT => \N__6436\,
            PACKAGEPIN => cpureset_wire
        );

    \arse.io_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6438\,
            PADOUT => \N__6437\,
            PADIN => \N__6436\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5579\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5915\
        );

    \lcol3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6429\,
            DIN => \N__6428\,
            DOUT => \N__6427\,
            PACKAGEPIN => lcol3_wire
        );

    \lcol3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6429\,
            PADOUT => \N__6428\,
            PADIN => \N__6427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2555\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \deldn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6420\,
            DIN => \N__6419\,
            DOUT => \N__6418\,
            PACKAGEPIN => deldn_wire
        );

    \deldn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6420\,
            PADOUT => \N__6419\,
            PADIN => \N__6418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => deldn_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6411\,
            DIN => \N__6410\,
            DOUT => \N__6409\,
            PACKAGEPIN => led2_wire
        );

    \led2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6411\,
            PADOUT => \N__6410\,
            PADIN => \N__6409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4811\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delup_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6402\,
            DIN => \N__6401\,
            DOUT => \N__6400\,
            PACKAGEPIN => delup_wire
        );

    \delup_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6402\,
            PADOUT => \N__6401\,
            PADIN => \N__6400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delup_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led6_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6393\,
            DIN => \N__6392\,
            DOUT => \N__6391\,
            PACKAGEPIN => led6_wire
        );

    \led6_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6393\,
            PADOUT => \N__6392\,
            PADIN => \N__6391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3668\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led8_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6384\,
            DIN => \N__6383\,
            DOUT => \N__6382\,
            PACKAGEPIN => led8_wire
        );

    \led8_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6384\,
            PADOUT => \N__6383\,
            PADIN => \N__6382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3626\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6375\,
            DIN => \N__6374\,
            DOUT => \N__6373\,
            PACKAGEPIN => led4_wire
        );

    \led4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6375\,
            PADOUT => \N__6374\,
            PADIN => \N__6373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6366\,
            DIN => \N__6365\,
            DOUT => \N__6364\,
            PACKAGEPIN => apureset_wire
        );

    \arse.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6366\,
            PADOUT => \N__6365\,
            PADIN => \N__6364\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6080\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5914\
        );

    \lcol4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6357\,
            DIN => \N__6356\,
            DOUT => \N__6355\,
            PACKAGEPIN => lcol4_wire
        );

    \lcol4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6357\,
            PADOUT => \N__6356\,
            PADIN => \N__6355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2540\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.diveight.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6348\,
            DIN => \N__6347\,
            DOUT => \N__6346\,
            PACKAGEPIN => cpuclk_wire
        );

    \arse.diveight.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6348\,
            PADOUT => \N__6347\,
            PADIN => \N__6346\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__5975\,
            OUTPUTENABLE => \N__4972\,
            DIN0 => OPEN,
            DOUT0 => \N__5804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5914\
        );

    \led5_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6339\,
            DIN => \N__6338\,
            DOUT => \N__6337\,
            PACKAGEPIN => led5_wire
        );

    \led5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6339\,
            PADOUT => \N__6338\,
            PADIN => \N__6337\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4968\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \consolereset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6330\,
            DIN => \N__6329\,
            DOUT => \N__6328\,
            PACKAGEPIN => consolereset_wire
        );

    \consolereset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6330\,
            PADOUT => \N__6329\,
            PADIN => \N__6328\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => consolereset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6321\,
            DIN => \N__6320\,
            DOUT => \N__6319\,
            PACKAGEPIN => lcol2_wire
        );

    \lcol2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6321\,
            PADOUT => \N__6320\,
            PADIN => \N__6319\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3341\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6312\,
            DIN => \N__6311\,
            DOUT => \N__6310\,
            PACKAGEPIN => led1_wire
        );

    \led1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6312\,
            PADOUT => \N__6311\,
            PADIN => \N__6310\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4949\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \apusync_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6303\,
            DIN => \N__6302\,
            DOUT => \N__6301\,
            PACKAGEPIN => apusync_wire
        );

    \apusync_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6303\,
            PADOUT => \N__6302\,
            PADIN => \N__6301\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => apusync_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6294\,
            DIN => \N__6293\,
            DOUT => \N__6292\,
            PACKAGEPIN => led7_wire
        );

    \led7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6294\,
            PADOUT => \N__6293\,
            PADIN => \N__6292\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3758\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6285\,
            DIN => \N__6284\,
            DOUT => \N__6283\,
            PACKAGEPIN => lcol1_wire
        );

    \lcol1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6285\,
            PADOUT => \N__6284\,
            PADIN => \N__6283\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__6266\,
            I => \N__6261\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__6265\,
            I => \N__6258\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6252\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6245\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6245\
        );

    \I__1500\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6245\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6240\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6240\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6252\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6245\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6240\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__6233\,
            I => \N__6226\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6222\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6211\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6211\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6211\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6211\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6211\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6222\,
            I => \arse.divseven.sevenZ0\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6211\,
            I => \arse.divseven.sevenZ0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1483\ : Span12Mux_v
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__1482\ : Odrv12
    port map (
            O => \N__6197\,
            I => apusync_c
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6186\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6183\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6180\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6186\,
            I => \N__6175\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6183\,
            I => \N__6170\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6180\,
            I => \N__6170\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6167\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6164\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__6175\,
            I => \N__6157\
        );

    \I__1471\ : Span4Mux_h
    port map (
            O => \N__6170\,
            I => \N__6157\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6157\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6164\,
            I => \N__6154\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__6157\,
            I => \N__6148\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__6154\,
            I => \N__6148\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6145\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__6148\,
            I => \arse.apusynclatchedZ0\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6145\,
            I => \arse.apusynclatchedZ0\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__1461\ : Span4Mux_v
    port map (
            O => \N__6134\,
            I => \N__6129\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6126\
        );

    \I__1459\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6123\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__6129\,
            I => \N__6120\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6126\,
            I => \N__6117\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6123\,
            I => \N__6114\
        );

    \I__1455\ : Sp12to4
    port map (
            O => \N__6120\,
            I => \N__6111\
        );

    \I__1454\ : Span4Mux_v
    port map (
            O => \N__6117\,
            I => \N__6108\
        );

    \I__1453\ : Span12Mux_s10_h
    port map (
            O => \N__6114\,
            I => \N__6104\
        );

    \I__1452\ : Span12Mux_v
    port map (
            O => \N__6111\,
            I => \N__6099\
        );

    \I__1451\ : Sp12to4
    port map (
            O => \N__6108\,
            I => \N__6099\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__6107\,
            I => \N__6096\
        );

    \I__1449\ : Span12Mux_v
    port map (
            O => \N__6104\,
            I => \N__6093\
        );

    \I__1448\ : Span12Mux_h
    port map (
            O => \N__6099\,
            I => \N__6090\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6087\
        );

    \I__1446\ : Odrv12
    port map (
            O => \N__6093\,
            I => debouncedconsolereset
        );

    \I__1445\ : Odrv12
    port map (
            O => \N__6090\,
            I => debouncedconsolereset
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6087\,
            I => debouncedconsolereset
        );

    \I__1443\ : IoInMux
    port map (
            O => \N__6080\,
            I => \N__6077\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6077\,
            I => \arse.apuresetoutregZ0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6070\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__6073\,
            I => \N__6067\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6062\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6055\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6055\
        );

    \I__1436\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6055\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__6062\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6055\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6045\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6042\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6036\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6045\,
            I => \N__6031\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6042\,
            I => \N__6031\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6024\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6024\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6024\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6036\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1424\ : Odrv12
    port map (
            O => \N__6031\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6024\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6011\,
            I => \N__6006\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6010\,
            I => \N__6001\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6001\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__6006\,
            I => \arse.diveight.counterZ0Z_1\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6001\,
            I => \arse.diveight.counterZ0Z_1\
        );

    \I__1415\ : InMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5988\
        );

    \I__1413\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5985\
        );

    \I__1412\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5982\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__5988\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__5985\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__5982\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__1408\ : IoInMux
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__5972\,
            I => \arse.diveight.doutZ0Z_1\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1405\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__5963\,
            I => \arse.divseven.N_46_0\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__5960\,
            I => \N__5955\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__5959\,
            I => \N__5949\
        );

    \I__1401\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5946\
        );

    \I__1400\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5939\
        );

    \I__1399\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5939\
        );

    \I__1398\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5939\
        );

    \I__1397\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5934\
        );

    \I__1396\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5934\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__5946\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__5939\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__5934\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1392\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5923\
        );

    \I__1391\ : IoInMux
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__5923\,
            I => \arse.divseven.doutZ0Z_1\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__5920\,
            I => \arse.divseven.doutZ0Z_1\
        );

    \I__1388\ : ClkMux
    port map (
            O => \N__5915\,
            I => \N__5870\
        );

    \I__1387\ : ClkMux
    port map (
            O => \N__5914\,
            I => \N__5870\
        );

    \I__1386\ : ClkMux
    port map (
            O => \N__5913\,
            I => \N__5870\
        );

    \I__1385\ : ClkMux
    port map (
            O => \N__5912\,
            I => \N__5870\
        );

    \I__1384\ : ClkMux
    port map (
            O => \N__5911\,
            I => \N__5870\
        );

    \I__1383\ : ClkMux
    port map (
            O => \N__5910\,
            I => \N__5870\
        );

    \I__1382\ : ClkMux
    port map (
            O => \N__5909\,
            I => \N__5870\
        );

    \I__1381\ : ClkMux
    port map (
            O => \N__5908\,
            I => \N__5870\
        );

    \I__1380\ : ClkMux
    port map (
            O => \N__5907\,
            I => \N__5870\
        );

    \I__1379\ : ClkMux
    port map (
            O => \N__5906\,
            I => \N__5870\
        );

    \I__1378\ : ClkMux
    port map (
            O => \N__5905\,
            I => \N__5870\
        );

    \I__1377\ : ClkMux
    port map (
            O => \N__5904\,
            I => \N__5870\
        );

    \I__1376\ : ClkMux
    port map (
            O => \N__5903\,
            I => \N__5870\
        );

    \I__1375\ : ClkMux
    port map (
            O => \N__5902\,
            I => \N__5870\
        );

    \I__1374\ : ClkMux
    port map (
            O => \N__5901\,
            I => \N__5870\
        );

    \I__1373\ : GlobalMux
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__1372\ : gio2CtrlBuf
    port map (
            O => \N__5867\,
            I => \PLLOUTCORE_g\
        );

    \I__1371\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5855\
        );

    \I__1370\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5852\
        );

    \I__1369\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5841\
        );

    \I__1368\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5841\
        );

    \I__1367\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5841\
        );

    \I__1366\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5841\
        );

    \I__1365\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5841\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__5855\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5852\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__5841\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1361\ : IoInMux
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__5831\,
            I => \arse.divseven.doutZ0Z_0\
        );

    \I__1359\ : CEMux
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__5822\,
            I => \arse.divseven.un1_dout_2_sqmuxa_0_i\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__5819\,
            I => \N__5815\
        );

    \I__1355\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5812\
        );

    \I__1354\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5809\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5812\,
            I => \arse.doingsevenZ0\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__5809\,
            I => \arse.doingsevenZ0\
        );

    \I__1351\ : IoInMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__1349\ : Span4Mux_s0_h
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__5795\,
            I => \arse.diveight.doutZ1Z_0\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__5789\,
            I => \arse.divseven.un1_counter_i_0_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5781\
        );

    \I__1344\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5776\
        );

    \I__1343\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5773\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__5781\,
            I => \N__5770\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5765\
        );

    \I__1340\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5765\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5760\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__5773\,
            I => \N__5760\
        );

    \I__1337\ : Span4Mux_h
    port map (
            O => \N__5770\,
            I => \N__5756\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__5765\,
            I => \N__5751\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__5760\,
            I => \N__5751\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5748\
        );

    \I__1333\ : Span4Mux_h
    port map (
            O => \N__5756\,
            I => \N__5745\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__5751\,
            I => \delayConstantZ0Z_4\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__5748\,
            I => \delayConstantZ0Z_4\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__5745\,
            I => \delayConstantZ0Z_4\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5734\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__5737\,
            I => \N__5730\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5734\,
            I => \N__5725\
        );

    \I__1326\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5722\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5719\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5716\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5713\
        );

    \I__1322\ : Span4Mux_v
    port map (
            O => \N__5725\,
            I => \N__5709\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__5722\,
            I => \N__5705\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__5719\,
            I => \N__5698\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N__5698\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5698\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5694\
        );

    \I__1316\ : Sp12to4
    port map (
            O => \N__5709\,
            I => \N__5691\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5688\
        );

    \I__1314\ : Span4Mux_v
    port map (
            O => \N__5705\,
            I => \N__5683\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__5698\,
            I => \N__5683\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5680\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5694\,
            I => \delayConstantZ0Z_0\
        );

    \I__1310\ : Odrv12
    port map (
            O => \N__5691\,
            I => \delayConstantZ0Z_0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5688\,
            I => \delayConstantZ0Z_0\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__5683\,
            I => \delayConstantZ0Z_0\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5680\,
            I => \delayConstantZ0Z_0\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5663\,
            I => \N__5657\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5654\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5651\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5648\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__5657\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5654\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__5651\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5648\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__5639\,
            I => \N__5633\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5630\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5627\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5624\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5621\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5630\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5627\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5624\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5621\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5609\,
            I => \arse.g0_3\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__5606\,
            I => \arse.g0_2_cascade_\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5600\,
            I => \arse.g0_4\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5594\,
            I => \arse.N_6\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5588\,
            I => \arse.g0_1\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__5585\,
            I => \arse.g0_7_cascade_\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__5582\,
            I => \arse.cpuresetoutreg_1_sqmuxa_cascade_\
        );

    \I__1276\ : IoInMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5576\,
            I => \N__5572\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5569\
        );

    \I__1273\ : Span4Mux_s3_h
    port map (
            O => \N__5572\,
            I => \N__5566\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5569\,
            I => \arse.cpuresetoutregZ0\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__5566\,
            I => \arse.cpuresetoutregZ0\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5558\,
            I => \arse.doingseven4\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5552\,
            I => \arse.doingseven3\
        );

    \I__1266\ : SRMux
    port map (
            O => \N__5549\,
            I => \N__5544\
        );

    \I__1265\ : SRMux
    port map (
            O => \N__5548\,
            I => \N__5541\
        );

    \I__1264\ : SRMux
    port map (
            O => \N__5547\,
            I => \N__5537\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5544\,
            I => \N__5534\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5541\,
            I => \N__5531\
        );

    \I__1261\ : SRMux
    port map (
            O => \N__5540\,
            I => \N__5528\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5525\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__5534\,
            I => debouncedconsolereset_i
        );

    \I__1258\ : Odrv12
    port map (
            O => \N__5531\,
            I => debouncedconsolereset_i
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5528\,
            I => debouncedconsolereset_i
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__5525\,
            I => debouncedconsolereset_i
        );

    \I__1255\ : InMux
    port map (
            O => \N__5516\,
            I => \arse.un1_cpuresetcount_1_cry_6\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__5513\,
            I => \N__5509\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__5512\,
            I => \N__5503\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5497\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5497\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5490\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5486\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5481\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5481\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5478\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5473\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5473\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__5494\,
            I => \N__5470\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__5493\,
            I => \N__5467\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5463\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5460\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5486\,
            I => \N__5457\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5481\,
            I => \N__5450\
        );

    \I__1237\ : Span4Mux_h
    port map (
            O => \N__5478\,
            I => \N__5450\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5450\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5447\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5442\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5442\
        );

    \I__1232\ : Span12Mux_s11_h
    port map (
            O => \N__5463\,
            I => \N__5437\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5460\,
            I => \N__5437\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__5457\,
            I => \N__5432\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__5450\,
            I => \N__5432\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5447\,
            I => \delayConstantZ0Z_1\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__5442\,
            I => \delayConstantZ0Z_1\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__5437\,
            I => \delayConstantZ0Z_1\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__5432\,
            I => \delayConstantZ0Z_1\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5411\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__5419\,
            I => \N__5408\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__5418\,
            I => \N__5402\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__5417\,
            I => \N__5399\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__5416\,
            I => \N__5396\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__5415\,
            I => \N__5393\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__5414\,
            I => \N__5390\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5411\,
            I => \N__5387\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5382\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \N__5379\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__5406\,
            I => \N__5376\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5371\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5371\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5366\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5366\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5361\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5361\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__5387\,
            I => \N__5358\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5386\,
            I => \N__5355\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5352\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5382\,
            I => \N__5349\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5344\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5344\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5371\,
            I => \N__5337\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5337\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5361\,
            I => \N__5337\
        );

    \I__1197\ : Sp12to4
    port map (
            O => \N__5358\,
            I => \N__5334\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5331\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5352\,
            I => \N__5322\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__5349\,
            I => \N__5322\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5322\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__5337\,
            I => \N__5322\
        );

    \I__1191\ : Odrv12
    port map (
            O => \N__5334\,
            I => \delayConstantZ0Z_5\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5331\,
            I => \delayConstantZ0Z_5\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__5322\,
            I => \delayConstantZ0Z_5\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5312\,
            I => \arse.g0_i_a3_4\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5303\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5300\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5297\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5294\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5303\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5300\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5297\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5294\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__5285\,
            I => \arse.doingseven3_6_cascade_\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5276\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5273\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5270\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5267\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5276\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5273\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5270\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5267\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5255\,
            I => \arse.doingseven3_1\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5249\,
            I => \arse.doingseven3_6\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__5246\,
            I => \arse.doingseven3_1_cascade_\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__1161\ : Span4Mux_h
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__5231\,
            I => \delayConstant_fastZ0Z_6\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__1156\ : Span4Mux_h
    port map (
            O => \N__5219\,
            I => \N__5216\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__5216\,
            I => \delayConstant_fastZ0Z_2\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__5213\,
            I => \N__5207\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__5212\,
            I => \N__5204\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__5211\,
            I => \N__5201\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5198\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5195\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5190\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5190\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5198\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5195\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5190\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5175\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5175\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5172\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5169\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5175\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5172\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5169\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5159\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5159\,
            I => \N__5155\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__5158\,
            I => \N__5148\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__5155\,
            I => \N__5144\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5141\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__5153\,
            I => \N__5138\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5135\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5132\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5129\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5126\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__5144\,
            I => \N__5123\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5120\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5117\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5135\,
            I => \N__5112\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5132\,
            I => \N__5112\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5129\,
            I => \N__5107\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5126\,
            I => \N__5107\
        );

    \I__1120\ : Span4Mux_h
    port map (
            O => \N__5123\,
            I => \N__5102\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__5120\,
            I => \N__5102\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5117\,
            I => \delayConstantZ0Z_7\
        );

    \I__1117\ : Odrv12
    port map (
            O => \N__5112\,
            I => \delayConstantZ0Z_7\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__5107\,
            I => \delayConstantZ0Z_7\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__5102\,
            I => \delayConstantZ0Z_7\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5089\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__5092\,
            I => \N__5084\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5089\,
            I => \N__5079\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5076\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5073\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5070\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5065\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5065\
        );

    \I__1106\ : Span4Mux_h
    port map (
            O => \N__5079\,
            I => \N__5062\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5076\,
            I => \N__5059\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5073\,
            I => \N__5055\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5070\,
            I => \N__5052\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5049\
        );

    \I__1101\ : Span4Mux_v
    port map (
            O => \N__5062\,
            I => \N__5046\
        );

    \I__1100\ : Span4Mux_h
    port map (
            O => \N__5059\,
            I => \N__5043\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5040\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__5055\,
            I => \N__5037\
        );

    \I__1097\ : Span4Mux_v
    port map (
            O => \N__5052\,
            I => \N__5032\
        );

    \I__1096\ : Span4Mux_v
    port map (
            O => \N__5049\,
            I => \N__5032\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__5046\,
            I => \delayConstantZ0Z_3\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__5043\,
            I => \delayConstantZ0Z_3\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5040\,
            I => \delayConstantZ0Z_3\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__5037\,
            I => \delayConstantZ0Z_3\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__5032\,
            I => \delayConstantZ0Z_3\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__5021\,
            I => \N__5017\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5012\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5009\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5004\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5004\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5012\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5009\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5004\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4990\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4983\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4983\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4983\
        );

    \I__1078\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4980\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4990\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__4983\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4980\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1074\ : IoInMux
    port map (
            O => \N__4973\,
            I => \N__4969\
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__4972\,
            I => \N__4965\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4969\,
            I => \N__4962\
        );

    \I__1071\ : IoInMux
    port map (
            O => \N__4968\,
            I => \N__4959\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4965\,
            I => \N__4956\
        );

    \I__1069\ : Span4Mux_s3_h
    port map (
            O => \N__4962\,
            I => \N__4953\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__4959\,
            I => \N__4950\
        );

    \I__1067\ : IoSpan4Mux
    port map (
            O => \N__4956\,
            I => \N__4946\
        );

    \I__1066\ : Span4Mux_v
    port map (
            O => \N__4953\,
            I => \N__4943\
        );

    \I__1065\ : IoSpan4Mux
    port map (
            O => \N__4950\,
            I => \N__4940\
        );

    \I__1064\ : IoInMux
    port map (
            O => \N__4949\,
            I => \N__4937\
        );

    \I__1063\ : Sp12to4
    port map (
            O => \N__4946\,
            I => \N__4934\
        );

    \I__1062\ : Sp12to4
    port map (
            O => \N__4943\,
            I => \N__4931\
        );

    \I__1061\ : IoSpan4Mux
    port map (
            O => \N__4940\,
            I => \N__4928\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4937\,
            I => \N__4925\
        );

    \I__1059\ : Span12Mux_s9_h
    port map (
            O => \N__4934\,
            I => \N__4922\
        );

    \I__1058\ : Span12Mux_s9_h
    port map (
            O => \N__4931\,
            I => \N__4919\
        );

    \I__1057\ : Span4Mux_s1_v
    port map (
            O => \N__4928\,
            I => \N__4914\
        );

    \I__1056\ : Span4Mux_s1_v
    port map (
            O => \N__4925\,
            I => \N__4914\
        );

    \I__1055\ : Span12Mux_v
    port map (
            O => \N__4922\,
            I => \N__4911\
        );

    \I__1054\ : Span12Mux_v
    port map (
            O => \N__4919\,
            I => \N__4908\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__4914\,
            I => \N__4905\
        );

    \I__1052\ : Odrv12
    port map (
            O => \N__4911\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1051\ : Odrv12
    port map (
            O => \N__4908\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1050\ : Odrv4
    port map (
            O => \N__4905\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4898\,
            I => \arse.un1_cpuresetcount_1_cry_0\
        );

    \I__1048\ : InMux
    port map (
            O => \N__4895\,
            I => \arse.un1_cpuresetcount_1_cry_1\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4892\,
            I => \arse.un1_cpuresetcount_1_cry_2\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4889\,
            I => \arse.un1_cpuresetcount_1_cry_3\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4886\,
            I => \arse.un1_cpuresetcount_1_cry_4\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4883\,
            I => \arse.un1_cpuresetcount_1_cry_5\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4877\,
            I => \dig1.N_25\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__4874\,
            I => \dig1.N_22_cascade_\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4868\,
            I => \dig1.leds_17_i_0_ns_1_2\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4861\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4858\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4861\,
            I => \un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4858\,
            I => \un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4849\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4846\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4849\,
            I => \un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4846\,
            I => \un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92\
        );

    \I__1030\ : SRMux
    port map (
            O => \N__4841\,
            I => \N__4817\
        );

    \I__1029\ : SRMux
    port map (
            O => \N__4840\,
            I => \N__4817\
        );

    \I__1028\ : SRMux
    port map (
            O => \N__4839\,
            I => \N__4817\
        );

    \I__1027\ : SRMux
    port map (
            O => \N__4838\,
            I => \N__4817\
        );

    \I__1026\ : SRMux
    port map (
            O => \N__4837\,
            I => \N__4817\
        );

    \I__1025\ : SRMux
    port map (
            O => \N__4836\,
            I => \N__4817\
        );

    \I__1024\ : SRMux
    port map (
            O => \N__4835\,
            I => \N__4817\
        );

    \I__1023\ : SRMux
    port map (
            O => \N__4834\,
            I => \N__4817\
        );

    \I__1022\ : GlobalMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__1021\ : gio2CtrlBuf
    port map (
            O => \N__4814\,
            I => masterreset_c_i_g
        );

    \I__1020\ : IoInMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__1018\ : IoSpan4Mux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__1017\ : Span4Mux_s3_v
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__1016\ : Sp12to4
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__1015\ : Span12Mux_s11_v
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__1014\ : Odrv12
    port map (
            O => \N__4793\,
            I => leds_1_i_0_1
        );

    \I__1013\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4787\,
            I => \N__4757\
        );

    \I__1011\ : ClkMux
    port map (
            O => \N__4786\,
            I => \N__4700\
        );

    \I__1010\ : ClkMux
    port map (
            O => \N__4785\,
            I => \N__4700\
        );

    \I__1009\ : ClkMux
    port map (
            O => \N__4784\,
            I => \N__4700\
        );

    \I__1008\ : ClkMux
    port map (
            O => \N__4783\,
            I => \N__4700\
        );

    \I__1007\ : ClkMux
    port map (
            O => \N__4782\,
            I => \N__4700\
        );

    \I__1006\ : ClkMux
    port map (
            O => \N__4781\,
            I => \N__4700\
        );

    \I__1005\ : ClkMux
    port map (
            O => \N__4780\,
            I => \N__4700\
        );

    \I__1004\ : ClkMux
    port map (
            O => \N__4779\,
            I => \N__4700\
        );

    \I__1003\ : ClkMux
    port map (
            O => \N__4778\,
            I => \N__4700\
        );

    \I__1002\ : ClkMux
    port map (
            O => \N__4777\,
            I => \N__4700\
        );

    \I__1001\ : ClkMux
    port map (
            O => \N__4776\,
            I => \N__4700\
        );

    \I__1000\ : ClkMux
    port map (
            O => \N__4775\,
            I => \N__4700\
        );

    \I__999\ : ClkMux
    port map (
            O => \N__4774\,
            I => \N__4700\
        );

    \I__998\ : ClkMux
    port map (
            O => \N__4773\,
            I => \N__4700\
        );

    \I__997\ : ClkMux
    port map (
            O => \N__4772\,
            I => \N__4700\
        );

    \I__996\ : ClkMux
    port map (
            O => \N__4771\,
            I => \N__4700\
        );

    \I__995\ : ClkMux
    port map (
            O => \N__4770\,
            I => \N__4700\
        );

    \I__994\ : ClkMux
    port map (
            O => \N__4769\,
            I => \N__4700\
        );

    \I__993\ : ClkMux
    port map (
            O => \N__4768\,
            I => \N__4700\
        );

    \I__992\ : ClkMux
    port map (
            O => \N__4767\,
            I => \N__4700\
        );

    \I__991\ : ClkMux
    port map (
            O => \N__4766\,
            I => \N__4700\
        );

    \I__990\ : ClkMux
    port map (
            O => \N__4765\,
            I => \N__4700\
        );

    \I__989\ : ClkMux
    port map (
            O => \N__4764\,
            I => \N__4700\
        );

    \I__988\ : ClkMux
    port map (
            O => \N__4763\,
            I => \N__4700\
        );

    \I__987\ : ClkMux
    port map (
            O => \N__4762\,
            I => \N__4700\
        );

    \I__986\ : ClkMux
    port map (
            O => \N__4761\,
            I => \N__4700\
        );

    \I__985\ : ClkMux
    port map (
            O => \N__4760\,
            I => \N__4700\
        );

    \I__984\ : Glb2LocalMux
    port map (
            O => \N__4757\,
            I => \N__4700\
        );

    \I__983\ : GlobalMux
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__982\ : gio2CtrlBuf
    port map (
            O => \N__4697\,
            I => \PACKAGEPIN_0_c_g\
        );

    \I__981\ : CEMux
    port map (
            O => \N__4694\,
            I => \N__4691\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4691\,
            I => \N__4686\
        );

    \I__979\ : CEMux
    port map (
            O => \N__4690\,
            I => \N__4683\
        );

    \I__978\ : CEMux
    port map (
            O => \N__4689\,
            I => \N__4675\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__4686\,
            I => \N__4670\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4683\,
            I => \N__4670\
        );

    \I__975\ : CEMux
    port map (
            O => \N__4682\,
            I => \N__4667\
        );

    \I__974\ : CEMux
    port map (
            O => \N__4681\,
            I => \N__4657\
        );

    \I__973\ : CEMux
    port map (
            O => \N__4680\,
            I => \N__4654\
        );

    \I__972\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4651\
        );

    \I__971\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4648\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4675\,
            I => \N__4645\
        );

    \I__969\ : Span4Mux_h
    port map (
            O => \N__4670\,
            I => \N__4640\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4640\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \N__4634\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__4665\,
            I => \N__4630\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__4664\,
            I => \N__4626\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__4663\,
            I => \N__4623\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \N__4620\
        );

    \I__962\ : CEMux
    port map (
            O => \N__4661\,
            I => \N__4614\
        );

    \I__961\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4611\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4657\,
            I => \N__4606\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4654\,
            I => \N__4606\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4601\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4648\,
            I => \N__4601\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__4645\,
            I => \N__4596\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__4640\,
            I => \N__4596\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__4639\,
            I => \N__4592\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__4638\,
            I => \N__4589\
        );

    \I__952\ : InMux
    port map (
            O => \N__4637\,
            I => \N__4583\
        );

    \I__951\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4580\
        );

    \I__950\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4577\
        );

    \I__949\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4572\
        );

    \I__948\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4572\
        );

    \I__947\ : InMux
    port map (
            O => \N__4626\,
            I => \N__4569\
        );

    \I__946\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4564\
        );

    \I__945\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4564\
        );

    \I__944\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4557\
        );

    \I__943\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4557\
        );

    \I__942\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4557\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4554\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4611\,
            I => \N__4549\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__4606\,
            I => \N__4549\
        );

    \I__938\ : Span4Mux_h
    port map (
            O => \N__4601\,
            I => \N__4544\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__4596\,
            I => \N__4544\
        );

    \I__936\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4539\
        );

    \I__935\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4539\
        );

    \I__934\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4530\
        );

    \I__933\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4530\
        );

    \I__932\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4530\
        );

    \I__931\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4530\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4583\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4580\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4577\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4572\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4569\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4564\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4557\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__923\ : Odrv12
    port map (
            O => \N__4554\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4549\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__4544\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4539\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4530\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__4505\,
            I => \dig1.N_52_cascade_\
        );

    \I__917\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4499\,
            I => \dig1.N_54\
        );

    \I__915\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4493\,
            I => \dig1.N_55\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__4490\,
            I => \N__4485\
        );

    \I__912\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4480\
        );

    \I__911\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4480\
        );

    \I__910\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4477\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4467\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4460\
        );

    \I__907\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4455\
        );

    \I__906\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4455\
        );

    \I__905\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4440\
        );

    \I__904\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4435\
        );

    \I__903\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4435\
        );

    \I__902\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4432\
        );

    \I__901\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4429\
        );

    \I__900\ : Span4Mux_h
    port map (
            O => \N__4467\,
            I => \N__4426\
        );

    \I__899\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4421\
        );

    \I__898\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4421\
        );

    \I__897\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4416\
        );

    \I__896\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4416\
        );

    \I__895\ : Span4Mux_v
    port map (
            O => \N__4460\,
            I => \N__4411\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4455\,
            I => \N__4411\
        );

    \I__893\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4406\
        );

    \I__892\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4406\
        );

    \I__891\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4401\
        );

    \I__890\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4401\
        );

    \I__889\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4394\
        );

    \I__888\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4394\
        );

    \I__887\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4394\
        );

    \I__886\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4389\
        );

    \I__885\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4389\
        );

    \I__884\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4382\
        );

    \I__883\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4382\
        );

    \I__882\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4382\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4377\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4435\,
            I => \N__4377\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4432\,
            I => \colZ0Z_0\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4429\,
            I => \colZ0Z_0\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__4426\,
            I => \colZ0Z_0\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4421\,
            I => \colZ0Z_0\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4416\,
            I => \colZ0Z_0\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4411\,
            I => \colZ0Z_0\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4406\,
            I => \colZ0Z_0\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4401\,
            I => \colZ0Z_0\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4394\,
            I => \colZ0Z_0\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4389\,
            I => \colZ0Z_0\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4382\,
            I => \colZ0Z_0\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__4377\,
            I => \colZ0Z_0\
        );

    \I__867\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4344\
        );

    \I__866\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4344\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__4350\,
            I => \N__4341\
        );

    \I__864\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4338\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4344\,
            I => \N__4326\
        );

    \I__862\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4323\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4338\,
            I => \N__4319\
        );

    \I__860\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4314\
        );

    \I__859\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4314\
        );

    \I__858\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4301\
        );

    \I__857\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4296\
        );

    \I__856\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4296\
        );

    \I__855\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4291\
        );

    \I__854\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4291\
        );

    \I__853\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4288\
        );

    \I__852\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4285\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__4326\,
            I => \N__4282\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4323\,
            I => \N__4279\
        );

    \I__849\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4276\
        );

    \I__848\ : Span4Mux_v
    port map (
            O => \N__4319\,
            I => \N__4271\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4271\
        );

    \I__846\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4266\
        );

    \I__845\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4266\
        );

    \I__844\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4259\
        );

    \I__843\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4259\
        );

    \I__842\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4259\
        );

    \I__841\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4254\
        );

    \I__840\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4254\
        );

    \I__839\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4247\
        );

    \I__838\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4247\
        );

    \I__837\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4247\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4301\,
            I => \N__4240\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4296\,
            I => \N__4240\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4291\,
            I => \N__4240\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4288\,
            I => \colZ0Z_1\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4285\,
            I => \colZ0Z_1\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__4282\,
            I => \colZ0Z_1\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__4279\,
            I => \colZ0Z_1\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4276\,
            I => \colZ0Z_1\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__4271\,
            I => \colZ0Z_1\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4266\,
            I => \colZ0Z_1\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4259\,
            I => \colZ0Z_1\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4254\,
            I => \colZ0Z_1\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4247\,
            I => \colZ0Z_1\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__4240\,
            I => \colZ0Z_1\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4217\,
            I => \N__4209\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__4216\,
            I => \N__4205\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \N__4202\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__4214\,
            I => \N__4198\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4213\,
            I => \N__4192\
        );

    \I__817\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4187\
        );

    \I__816\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4187\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__4208\,
            I => \N__4184\
        );

    \I__814\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4179\
        );

    \I__813\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4179\
        );

    \I__812\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4176\
        );

    \I__811\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4173\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__4197\,
            I => \N__4169\
        );

    \I__809\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4166\
        );

    \I__808\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4161\
        );

    \I__807\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4161\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4187\,
            I => \N__4158\
        );

    \I__805\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4155\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4179\,
            I => \N__4152\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4176\,
            I => \N__4149\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4173\,
            I => \N__4146\
        );

    \I__801\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4141\
        );

    \I__800\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4141\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4166\,
            I => \N__4132\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4161\,
            I => \N__4132\
        );

    \I__797\ : Span4Mux_h
    port map (
            O => \N__4158\,
            I => \N__4132\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4155\,
            I => \N__4132\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__4152\,
            I => \N__4129\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__4149\,
            I => \delayConstantZ0Z_2\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__4146\,
            I => \delayConstantZ0Z_2\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4141\,
            I => \delayConstantZ0Z_2\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__4132\,
            I => \delayConstantZ0Z_2\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__4129\,
            I => \delayConstantZ0Z_2\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__4118\,
            I => \dig1.m47_ns_1_cascade_\
        );

    \I__788\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4108\
        );

    \I__787\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4105\
        );

    \I__786\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4102\
        );

    \I__785\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4099\
        );

    \I__784\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4096\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4108\,
            I => \N__4093\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4105\,
            I => col_1_1
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4102\,
            I => col_1_1
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4099\,
            I => col_1_1
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4096\,
            I => col_1_1
        );

    \I__778\ : Odrv4
    port map (
            O => \N__4093\,
            I => col_1_1
        );

    \I__777\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4079\,
            I => \dig1.N_49\
        );

    \I__775\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4073\,
            I => \dig1.m41_bm\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__4070\,
            I => \dig1.m41_am_cascade_\
        );

    \I__772\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4064\,
            I => \dig1.N_44\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__4061\,
            I => \dig1.m10_ns_1_cascade_\
        );

    \I__769\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4055\,
            I => \dig1.N_11_0\
        );

    \I__767\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4041\
        );

    \I__766\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4041\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4050\,
            I => \N__4033\
        );

    \I__764\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4028\
        );

    \I__763\ : InMux
    port map (
            O => \N__4048\,
            I => \N__4028\
        );

    \I__762\ : InMux
    port map (
            O => \N__4047\,
            I => \N__4023\
        );

    \I__761\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4023\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4041\,
            I => \N__4020\
        );

    \I__759\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4015\
        );

    \I__758\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4015\
        );

    \I__757\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4010\
        );

    \I__756\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4010\
        );

    \I__755\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4007\
        );

    \I__754\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4004\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4028\,
            I => \N__3999\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4023\,
            I => \N__3999\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__4020\,
            I => \N__3992\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4015\,
            I => \N__3992\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4010\,
            I => \N__3992\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4007\,
            I => \delayConstantZ0Z_6\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4004\,
            I => \delayConstantZ0Z_6\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__3999\,
            I => \delayConstantZ0Z_6\
        );

    \I__745\ : Odrv12
    port map (
            O => \N__3992\,
            I => \delayConstantZ0Z_6\
        );

    \I__744\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3980\,
            I => \olddn_RNIM5BH1Z0Z_1\
        );

    \I__742\ : InMux
    port map (
            O => \N__3977\,
            I => \un1_delayConstant_cry_0\
        );

    \I__741\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3971\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3971\,
            I => \olddn_RNIM5BHZ0Z1\
        );

    \I__739\ : InMux
    port map (
            O => \N__3968\,
            I => \un1_delayConstant_cry_1\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__3965\,
            I => \N__3962\
        );

    \I__737\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3959\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3959\,
            I => \olddn_RNIM5BH1Z0Z_2\
        );

    \I__735\ : InMux
    port map (
            O => \N__3956\,
            I => \un1_delayConstant_cry_2\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__733\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__3944\,
            I => \olddn_RNIM5BH1Z0Z_3\
        );

    \I__730\ : InMux
    port map (
            O => \N__3941\,
            I => \un1_delayConstant_cry_3\
        );

    \I__729\ : InMux
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3935\,
            I => \olddn_RNIM5BH1Z0Z_0\
        );

    \I__727\ : InMux
    port map (
            O => \N__3932\,
            I => \un1_delayConstant_cry_4\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__725\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3923\,
            I => \N__3920\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__3920\,
            I => \olddn_RNIM5BH1Z0Z_4\
        );

    \I__722\ : InMux
    port map (
            O => \N__3917\,
            I => \un1_delayConstant_cry_5\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__3914\,
            I => \N__3908\
        );

    \I__720\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3901\
        );

    \I__719\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3898\
        );

    \I__718\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3891\
        );

    \I__717\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3891\
        );

    \I__716\ : InMux
    port map (
            O => \N__3907\,
            I => \N__3891\
        );

    \I__715\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3884\
        );

    \I__714\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3884\
        );

    \I__713\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3884\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3901\,
            I => \delayConstant16_i\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3898\,
            I => \delayConstant16_i\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3891\,
            I => \delayConstant16_i\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3884\,
            I => \delayConstant16_i\
        );

    \I__708\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3864\
        );

    \I__707\ : InMux
    port map (
            O => \N__3874\,
            I => \N__3861\
        );

    \I__706\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3854\
        );

    \I__705\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3854\
        );

    \I__704\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3854\
        );

    \I__703\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3845\
        );

    \I__702\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3845\
        );

    \I__701\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3845\
        );

    \I__700\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3845\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3864\,
            I => \olddn_RNIEENHZ0\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3861\,
            I => \olddn_RNIEENHZ0\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3854\,
            I => \olddn_RNIEENHZ0\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3845\,
            I => \olddn_RNIEENHZ0\
        );

    \I__695\ : InMux
    port map (
            O => \N__3836\,
            I => \un1_delayConstant_cry_6\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__3833\,
            I => \dig1.N_15_cascade_\
        );

    \I__693\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3827\,
            I => \dig1.N_18\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__3824\,
            I => \N__3821\
        );

    \I__690\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3816\
        );

    \I__689\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3813\
        );

    \I__688\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3808\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3816\,
            I => \N__3803\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3813\,
            I => \N__3803\
        );

    \I__685\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3800\
        );

    \I__684\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3797\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3808\,
            I => slowclk
        );

    \I__682\ : Odrv4
    port map (
            O => \N__3803\,
            I => slowclk
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3800\,
            I => slowclk
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3797\,
            I => slowclk
        );

    \I__679\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3782\
        );

    \I__678\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3782\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3782\,
            I => \clock_out_RNIR6ER\
        );

    \I__676\ : InMux
    port map (
            O => \N__3779\,
            I => \N__3776\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3776\,
            I => \dig1.N_17\
        );

    \I__674\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3770\,
            I => \dig1.m32_bm\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__3767\,
            I => \N__3764\
        );

    \I__671\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3761\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3761\,
            I => \dig1.m32_am\
        );

    \I__669\ : IoInMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__667\ : Span4Mux_s2_v
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__666\ : Sp12to4
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__665\ : Span12Mux_h
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__664\ : Span12Mux_v
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__3740\,
            I => leds_1_i_2
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__661\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3731\,
            I => \un1_delayConstant_cry_0_c_RNOZ0\
        );

    \I__659\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3725\,
            I => \dig1.m77_am\
        );

    \I__657\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__655\ : Span4Mux_h
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3713\,
            I => \debounceup.out_cnv_2\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__652\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__650\ : Span12Mux_h
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__649\ : Span12Mux_v
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__3695\,
            I => delup_c
        );

    \I__647\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3687\
        );

    \I__646\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3682\
        );

    \I__645\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3682\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3687\,
            I => debouncedup
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3682\,
            I => debouncedup
        );

    \I__642\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__3671\,
            I => \dig1.m77_bm\
        );

    \I__639\ : IoInMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__637\ : IoSpan4Mux
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__636\ : IoSpan4Mux
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__635\ : Sp12to4
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__634\ : Span12Mux_s6_v
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__633\ : Odrv12
    port map (
            O => \N__3650\,
            I => leds_1_i_1
        );

    \I__632\ : IoInMux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__630\ : Span12Mux_s5_v
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__629\ : Span12Mux_v
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__3635\,
            I => lcol1_c
        );

    \I__627\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3629\,
            I => \dig1.N_39\
        );

    \I__625\ : IoInMux
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3623\,
            I => \N__3620\
        );

    \I__623\ : IoSpan4Mux
    port map (
            O => \N__3620\,
            I => \N__3617\
        );

    \I__622\ : Span4Mux_s3_v
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__621\ : Sp12to4
    port map (
            O => \N__3614\,
            I => \N__3611\
        );

    \I__620\ : Span12Mux_s10_v
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__619\ : Span12Mux_h
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__3605\,
            I => leds_1_i_3
        );

    \I__617\ : IoInMux
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__615\ : IoSpan4Mux
    port map (
            O => \N__3596\,
            I => \N__3592\
        );

    \I__614\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3589\
        );

    \I__613\ : Span4Mux_s2_v
    port map (
            O => \N__3592\,
            I => \N__3586\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3589\,
            I => \N__3580\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__3586\,
            I => \N__3577\
        );

    \I__610\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3574\
        );

    \I__609\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3571\
        );

    \I__608\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3568\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__3580\,
            I => \N__3565\
        );

    \I__606\ : Span4Mux_v
    port map (
            O => \N__3577\,
            I => \N__3560\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3574\,
            I => \N__3560\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3571\,
            I => \N__3554\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3568\,
            I => \N__3554\
        );

    \I__602\ : Span4Mux_h
    port map (
            O => \N__3565\,
            I => \N__3549\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__3560\,
            I => \N__3549\
        );

    \I__600\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3546\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__3554\,
            I => \N__3543\
        );

    \I__598\ : Sp12to4
    port map (
            O => \N__3549\,
            I => \N__3538\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3538\
        );

    \I__596\ : Sp12to4
    port map (
            O => \N__3543\,
            I => \N__3535\
        );

    \I__595\ : Span12Mux_h
    port map (
            O => \N__3538\,
            I => \N__3532\
        );

    \I__594\ : Span12Mux_h
    port map (
            O => \N__3535\,
            I => \N__3529\
        );

    \I__593\ : Span12Mux_v
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__592\ : Span12Mux_v
    port map (
            O => \N__3529\,
            I => \N__3523\
        );

    \I__591\ : Odrv12
    port map (
            O => \N__3526\,
            I => masterreset_c
        );

    \I__590\ : Odrv12
    port map (
            O => \N__3523\,
            I => masterreset_c
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3518\,
            I => \delayConstant16_i_cascade_\
        );

    \I__588\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3512\,
            I => \oldupZ0\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__585\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3501\
        );

    \I__584\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3496\
        );

    \I__583\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3496\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3501\,
            I => debounceddn
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3496\,
            I => debounceddn
        );

    \I__580\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3488\,
            I => \olddnZ0\
        );

    \I__578\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3482\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3482\,
            I => \dig1.N_72\
        );

    \I__576\ : InMux
    port map (
            O => \N__3479\,
            I => \N__3476\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__574\ : Span4Mux_h
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__3470\,
            I => \debouncedn.out_cnv_2\
        );

    \I__572\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__3461\,
            I => \N__3458\
        );

    \I__569\ : Sp12to4
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__568\ : Span12Mux_h
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__567\ : Span12Mux_v
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__3449\,
            I => deldn_c
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__3446\,
            I => \dig1.N_58_cascade_\
        );

    \I__564\ : InMux
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3440\,
            I => \dig1.leds_17_i_ns_1_2\
        );

    \I__562\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3434\,
            I => \dig1.N_61\
        );

    \I__560\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3428\,
            I => \dig1.m68_bm\
        );

    \I__558\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3422\,
            I => \dig1.m68_am\
        );

    \I__556\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3402\
        );

    \I__555\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3399\
        );

    \I__554\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3390\
        );

    \I__553\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3390\
        );

    \I__552\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3390\
        );

    \I__551\ : InMux
    port map (
            O => \N__3414\,
            I => \N__3381\
        );

    \I__550\ : InMux
    port map (
            O => \N__3413\,
            I => \N__3381\
        );

    \I__549\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3381\
        );

    \I__548\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3381\
        );

    \I__547\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3374\
        );

    \I__546\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3374\
        );

    \I__545\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3374\
        );

    \I__544\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3367\
        );

    \I__543\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3367\
        );

    \I__542\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3367\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3402\,
            I => \N__3362\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3399\,
            I => \N__3362\
        );

    \I__539\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3359\
        );

    \I__538\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3356\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3390\,
            I => \arses.counter8\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3381\,
            I => \arses.counter8\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3374\,
            I => \arses.counter8\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3367\,
            I => \arses.counter8\
        );

    \I__533\ : Odrv4
    port map (
            O => \N__3362\,
            I => \arses.counter8\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3359\,
            I => \arses.counter8\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3356\,
            I => \arses.counter8\
        );

    \I__530\ : IoInMux
    port map (
            O => \N__3341\,
            I => \N__3338\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3338\,
            I => \N__3335\
        );

    \I__528\ : IoSpan4Mux
    port map (
            O => \N__3335\,
            I => \N__3332\
        );

    \I__527\ : Span4Mux_s3_v
    port map (
            O => \N__3332\,
            I => \N__3329\
        );

    \I__526\ : Sp12to4
    port map (
            O => \N__3329\,
            I => \N__3326\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__524\ : Span12Mux_v
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__523\ : Odrv12
    port map (
            O => \N__3320\,
            I => lcol2_c
        );

    \I__522\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3313\
        );

    \I__521\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3310\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3313\,
            I => \arses.counterZ0Z_7\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3310\,
            I => \arses.counterZ0Z_7\
        );

    \I__518\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3301\
        );

    \I__517\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3298\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3301\,
            I => \arses.counterZ0Z_6\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3298\,
            I => \arses.counterZ0Z_6\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3293\,
            I => \N__3289\
        );

    \I__513\ : InMux
    port map (
            O => \N__3292\,
            I => \N__3286\
        );

    \I__512\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3283\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3286\,
            I => \arses.counterZ0Z_8\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3283\,
            I => \arses.counterZ0Z_8\
        );

    \I__509\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3274\
        );

    \I__508\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3271\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3274\,
            I => \arses.counterZ0Z_5\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3271\,
            I => \arses.counterZ0Z_5\
        );

    \I__505\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3262\
        );

    \I__504\ : InMux
    port map (
            O => \N__3265\,
            I => \N__3259\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3262\,
            I => \arses.counterZ0Z_4\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3259\,
            I => \arses.counterZ0Z_4\
        );

    \I__501\ : InMux
    port map (
            O => \N__3254\,
            I => \N__3249\
        );

    \I__500\ : InMux
    port map (
            O => \N__3253\,
            I => \N__3246\
        );

    \I__499\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3243\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3249\,
            I => \N__3240\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3246\,
            I => \N__3237\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3243\,
            I => \arses.counterZ0Z_1\
        );

    \I__495\ : Odrv4
    port map (
            O => \N__3240\,
            I => \arses.counterZ0Z_1\
        );

    \I__494\ : Odrv4
    port map (
            O => \N__3237\,
            I => \arses.counterZ0Z_1\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__3230\,
            I => \arses.un1_counterlto8_2_cascade_\
        );

    \I__492\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3223\
        );

    \I__491\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3220\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3223\,
            I => \arses.counterZ0Z_11\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3220\,
            I => \arses.counterZ0Z_11\
        );

    \I__488\ : InMux
    port map (
            O => \N__3215\,
            I => \N__3211\
        );

    \I__487\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3208\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3211\,
            I => \arses.counterZ0Z_10\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3208\,
            I => \arses.counterZ0Z_10\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__3203\,
            I => \arses.un1_counterlt11_cascade_\
        );

    \I__483\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3196\
        );

    \I__482\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3193\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3196\,
            I => \arses.counterZ0Z_9\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3193\,
            I => \arses.counterZ0Z_9\
        );

    \I__479\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3184\
        );

    \I__478\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3181\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3184\,
            I => \arses.counterZ0Z_14\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3181\,
            I => \arses.counterZ0Z_14\
        );

    \I__475\ : InMux
    port map (
            O => \N__3176\,
            I => \N__3172\
        );

    \I__474\ : InMux
    port map (
            O => \N__3175\,
            I => \N__3169\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3172\,
            I => \arses.counterZ0Z_13\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3169\,
            I => \arses.counterZ0Z_13\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__3164\,
            I => \arses.un1_counterlt13_0_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3157\
        );

    \I__469\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3157\,
            I => \arses.counterZ0Z_12\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3154\,
            I => \arses.counterZ0Z_12\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3149\,
            I => \arses.counter8_cascade_\
        );

    \I__465\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3142\
        );

    \I__464\ : InMux
    port map (
            O => \N__3145\,
            I => \N__3139\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3142\,
            I => \arses.counterZ0Z_3\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3139\,
            I => \arses.counterZ0Z_3\
        );

    \I__461\ : InMux
    port map (
            O => \N__3134\,
            I => \N__3130\
        );

    \I__460\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3127\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3130\,
            I => \arses.counterZ0Z_2\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3127\,
            I => \arses.counterZ0Z_2\
        );

    \I__457\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3119\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3119\,
            I => \arses.un1_counterlto4_2\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__454\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3108\
        );

    \I__453\ : InMux
    port map (
            O => \N__3112\,
            I => \N__3104\
        );

    \I__452\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3101\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3108\,
            I => \N__3098\
        );

    \I__450\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3095\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3104\,
            I => \arses.counterZ0Z_0\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3101\,
            I => \arses.counterZ0Z_0\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__3098\,
            I => \arses.counterZ0Z_0\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3095\,
            I => \arses.counterZ0Z_0\
        );

    \I__445\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3083\,
            I => \dig1.N_78\
        );

    \I__443\ : InMux
    port map (
            O => \N__3080\,
            I => \arses.un2_counter_cry_13\
        );

    \I__442\ : IoInMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__440\ : IoSpan4Mux
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__439\ : IoSpan4Mux
    port map (
            O => \N__3068\,
            I => \N__3065\
        );

    \I__438\ : Span4Mux_s3_v
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__437\ : Sp12to4
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__436\ : Span12Mux_s11_v
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__3056\,
            I => leds_1_i_0_3
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__3053\,
            I => \debounceup.counter_RNI45V02Z0Z_4_cascade_\
        );

    \I__433\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3042\
        );

    \I__432\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3042\
        );

    \I__431\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3039\
        );

    \I__430\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3036\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3042\,
            I => \debounceup.counterZ0Z_3\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3039\,
            I => \debounceup.counterZ0Z_3\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3036\,
            I => \debounceup.counterZ0Z_3\
        );

    \I__426\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3021\
        );

    \I__425\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3021\
        );

    \I__424\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3016\
        );

    \I__423\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3016\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3021\,
            I => \debounceup.counterZ0Z_2\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3016\,
            I => \debounceup.counterZ0Z_2\
        );

    \I__420\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3006\
        );

    \I__419\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3001\
        );

    \I__418\ : InMux
    port map (
            O => \N__3009\,
            I => \N__3001\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3006\,
            I => \debounceup.counterZ0Z_4\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3001\,
            I => \debounceup.counterZ0Z_4\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__2996\,
            I => \debounceup.counter18_0_2_cascade_\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2993\,
            I => \N__2989\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2992\,
            I => \N__2985\
        );

    \I__412\ : InMux
    port map (
            O => \N__2989\,
            I => \N__2981\
        );

    \I__411\ : InMux
    port map (
            O => \N__2988\,
            I => \N__2974\
        );

    \I__410\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2974\
        );

    \I__409\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2974\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2981\,
            I => \debounceup.counterZ0Z_0\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2974\,
            I => \debounceup.counterZ0Z_0\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__405\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2962\
        );

    \I__404\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2957\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2962\,
            I => \N__2954\
        );

    \I__402\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2949\
        );

    \I__401\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2949\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2957\,
            I => \debounceup.counter_RNI45V02Z0Z_4\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__2954\,
            I => \debounceup.counter_RNI45V02Z0Z_4\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2949\,
            I => \debounceup.counter_RNI45V02Z0Z_4\
        );

    \I__397\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2935\
        );

    \I__396\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2935\
        );

    \I__395\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2932\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2935\,
            I => \debounceup.counterZ0Z_1\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2932\,
            I => \debounceup.counterZ0Z_1\
        );

    \I__392\ : IoInMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__390\ : IoSpan4Mux
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__389\ : Span4Mux_s3_v
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__386\ : Span12Mux_v
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__2906\,
            I => leds_1_i_0_2
        );

    \I__384\ : InMux
    port map (
            O => \N__2903\,
            I => \arses.un2_counter_cry_3\
        );

    \I__383\ : InMux
    port map (
            O => \N__2900\,
            I => \arses.un2_counter_cry_4\
        );

    \I__382\ : InMux
    port map (
            O => \N__2897\,
            I => \arses.un2_counter_cry_5\
        );

    \I__381\ : InMux
    port map (
            O => \N__2894\,
            I => \arses.un2_counter_cry_6\
        );

    \I__380\ : InMux
    port map (
            O => \N__2891\,
            I => \arses.un2_counter_cry_7\
        );

    \I__379\ : InMux
    port map (
            O => \N__2888\,
            I => \bfn_17_17_0_\
        );

    \I__378\ : InMux
    port map (
            O => \N__2885\,
            I => \arses.un2_counter_cry_9\
        );

    \I__377\ : InMux
    port map (
            O => \N__2882\,
            I => \arses.un2_counter_cry_10\
        );

    \I__376\ : InMux
    port map (
            O => \N__2879\,
            I => \arses.un2_counter_cry_11\
        );

    \I__375\ : InMux
    port map (
            O => \N__2876\,
            I => \arses.un2_counter_cry_12\
        );

    \I__374\ : InMux
    port map (
            O => \N__2873\,
            I => \debounceconsolereset.un3_counter_cry_3\
        );

    \I__373\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2865\
        );

    \I__372\ : InMux
    port map (
            O => \N__2869\,
            I => \N__2860\
        );

    \I__371\ : InMux
    port map (
            O => \N__2868\,
            I => \N__2860\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2865\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2860\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__2855\,
            I => \clock_out_RNIR6ER_0_cascade_\
        );

    \I__367\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2849\,
            I => \debounceconsolereset.un3_counter_cry_2_THRU_CO\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2846\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__2843\,
            I => \N__2838\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__2842\,
            I => \N__2834\
        );

    \I__362\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2831\
        );

    \I__361\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2826\
        );

    \I__360\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2826\
        );

    \I__359\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2823\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2831\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2826\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2823\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__2816\,
            I => \N__2812\
        );

    \I__354\ : InMux
    port map (
            O => \N__2815\,
            I => \N__2807\
        );

    \I__353\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2804\
        );

    \I__352\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2799\
        );

    \I__351\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2799\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2807\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2804\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2799\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__346\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2786\,
            I => \debounceconsolereset.un3_counter_cry_1_THRU_CO\
        );

    \I__344\ : InMux
    port map (
            O => \N__2783\,
            I => \N__2777\
        );

    \I__343\ : InMux
    port map (
            O => \N__2782\,
            I => \N__2772\
        );

    \I__342\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2772\
        );

    \I__341\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2769\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2777\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2772\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2769\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__337\ : InMux
    port map (
            O => \N__2762\,
            I => \arses.un2_counter_cry_1\
        );

    \I__336\ : InMux
    port map (
            O => \N__2759\,
            I => \arses.un2_counter_cry_2\
        );

    \I__335\ : InMux
    port map (
            O => \N__2756\,
            I => \debounceup.un3_counter_cry_1\
        );

    \I__334\ : InMux
    port map (
            O => \N__2753\,
            I => \debounceup.un3_counter_cry_2\
        );

    \I__333\ : InMux
    port map (
            O => \N__2750\,
            I => \debounceup.un3_counter_cry_3\
        );

    \I__332\ : InMux
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2744\,
            I => \debounceup.un3_counter_cry_2_THRU_CO\
        );

    \I__330\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2738\,
            I => \debounceup.un3_counter_cry_1_THRU_CO\
        );

    \I__328\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2728\
        );

    \I__327\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2728\
        );

    \I__326\ : InMux
    port map (
            O => \N__2733\,
            I => \N__2725\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2728\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2725\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__2720\,
            I => \N__2716\
        );

    \I__322\ : CascadeMux
    port map (
            O => \N__2719\,
            I => \N__2711\
        );

    \I__321\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2704\
        );

    \I__320\ : InMux
    port map (
            O => \N__2715\,
            I => \N__2704\
        );

    \I__319\ : InMux
    port map (
            O => \N__2714\,
            I => \N__2704\
        );

    \I__318\ : InMux
    port map (
            O => \N__2711\,
            I => \N__2701\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2704\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2701\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__315\ : InMux
    port map (
            O => \N__2696\,
            I => \debounceconsolereset.un3_counter_cry_1\
        );

    \I__314\ : InMux
    port map (
            O => \N__2693\,
            I => \debounceconsolereset.un3_counter_cry_2\
        );

    \I__313\ : CascadeMux
    port map (
            O => \N__2690\,
            I => \debouncedn.counter_RNIBTPA2Z0Z_4_cascade_\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__2687\,
            I => \N__2681\
        );

    \I__311\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2678\
        );

    \I__310\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2673\
        );

    \I__309\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2673\
        );

    \I__308\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2670\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2678\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2673\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2670\,
            I => \debouncedn.counterZ0Z_0\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2663\,
            I => \debounceconsolereset.counter18_0_2_cascade_\
        );

    \I__303\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2657\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2657\,
            I => \debouncedn.un3_counter_cry_2_THRU_CO\
        );

    \I__301\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2648\
        );

    \I__300\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2643\
        );

    \I__299\ : InMux
    port map (
            O => \N__2652\,
            I => \N__2643\
        );

    \I__298\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2640\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2648\,
            I => \debouncedn.counterZ0Z_3\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2643\,
            I => \debouncedn.counterZ0Z_3\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2640\,
            I => \debouncedn.counterZ0Z_3\
        );

    \I__294\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2630\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2630\,
            I => \debouncedn.un3_counter_cry_1_THRU_CO\
        );

    \I__292\ : CascadeMux
    port map (
            O => \N__2627\,
            I => \N__2623\
        );

    \I__291\ : InMux
    port map (
            O => \N__2626\,
            I => \N__2618\
        );

    \I__290\ : InMux
    port map (
            O => \N__2623\,
            I => \N__2615\
        );

    \I__289\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2610\
        );

    \I__288\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2610\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2618\,
            I => \debouncedn.counter_RNIBTPA2Z0Z_4\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2615\,
            I => \debouncedn.counter_RNIBTPA2Z0Z_4\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2610\,
            I => \debouncedn.counter_RNIBTPA2Z0Z_4\
        );

    \I__284\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2595\
        );

    \I__283\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2595\
        );

    \I__282\ : InMux
    port map (
            O => \N__2601\,
            I => \N__2592\
        );

    \I__281\ : InMux
    port map (
            O => \N__2600\,
            I => \N__2589\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2595\,
            I => \debouncedn.counterZ0Z_2\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2592\,
            I => \debouncedn.counterZ0Z_2\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2589\,
            I => \debouncedn.counterZ0Z_2\
        );

    \I__277\ : InMux
    port map (
            O => \N__2582\,
            I => \N__2579\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__275\ : Span4Mux_v
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__274\ : Sp12to4
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__273\ : Span12Mux_h
    port map (
            O => \N__2570\,
            I => \N__2567\
        );

    \I__272\ : Span12Mux_v
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__271\ : Odrv12
    port map (
            O => \N__2564\,
            I => consolereset_c
        );

    \I__270\ : InMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2558\,
            I => \debounceconsolereset.out_cnv_2\
        );

    \I__268\ : IoInMux
    port map (
            O => \N__2555\,
            I => \N__2552\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__266\ : Sp12to4
    port map (
            O => \N__2549\,
            I => \N__2546\
        );

    \I__265\ : Span12Mux_s6_v
    port map (
            O => \N__2546\,
            I => \N__2543\
        );

    \I__264\ : Odrv12
    port map (
            O => \N__2543\,
            I => lcol3_c
        );

    \I__263\ : IoInMux
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__261\ : IoSpan4Mux
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__260\ : IoSpan4Mux
    port map (
            O => \N__2531\,
            I => \N__2528\
        );

    \I__259\ : Span4Mux_s3_v
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__258\ : Sp12to4
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__257\ : Odrv12
    port map (
            O => \N__2522\,
            I => lcol4_c
        );

    \I__256\ : InMux
    port map (
            O => \N__2519\,
            I => \debouncedn.un3_counter_cry_1\
        );

    \I__255\ : InMux
    port map (
            O => \N__2516\,
            I => \debouncedn.un3_counter_cry_2\
        );

    \I__254\ : InMux
    port map (
            O => \N__2513\,
            I => \debouncedn.un3_counter_cry_3\
        );

    \I__253\ : IoInMux
    port map (
            O => \N__2510\,
            I => \N__2507\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2507\,
            I => \N__2504\
        );

    \I__251\ : IoSpan4Mux
    port map (
            O => \N__2504\,
            I => \N__2501\
        );

    \I__250\ : Odrv4
    port map (
            O => \N__2501\,
            I => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__2498\,
            I => \debouncedn.counter18_0_2_cascade_\
        );

    \I__248\ : InMux
    port map (
            O => \N__2495\,
            I => \N__2490\
        );

    \I__247\ : InMux
    port map (
            O => \N__2494\,
            I => \N__2487\
        );

    \I__246\ : InMux
    port map (
            O => \N__2493\,
            I => \N__2484\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2490\,
            I => \debouncedn.counterZ0Z_1\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2487\,
            I => \debouncedn.counterZ0Z_1\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2484\,
            I => \debouncedn.counterZ0Z_1\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2477\,
            I => \N__2472\
        );

    \I__241\ : InMux
    port map (
            O => \N__2476\,
            I => \N__2469\
        );

    \I__240\ : InMux
    port map (
            O => \N__2475\,
            I => \N__2466\
        );

    \I__239\ : InMux
    port map (
            O => \N__2472\,
            I => \N__2463\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2469\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2466\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2463\,
            I => \debouncedn.counterZ0Z_4\
        );

    \I__235\ : IoInMux
    port map (
            O => \N__2456\,
            I => \N__2453\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2453\,
            I => \N__2450\
        );

    \I__233\ : IoSpan4Mux
    port map (
            O => \N__2450\,
            I => \N__2447\
        );

    \I__232\ : Span4Mux_s2_v
    port map (
            O => \N__2447\,
            I => \N__2444\
        );

    \I__231\ : Sp12to4
    port map (
            O => \N__2444\,
            I => \N__2441\
        );

    \I__230\ : Span12Mux_s10_v
    port map (
            O => \N__2441\,
            I => \N__2438\
        );

    \I__229\ : Span12Mux_v
    port map (
            O => \N__2438\,
            I => \N__2435\
        );

    \I__228\ : Span12Mux_h
    port map (
            O => \N__2435\,
            I => \N__2432\
        );

    \I__227\ : Odrv12
    port map (
            O => \N__2432\,
            I => \arse.divseven.io_0_D_IN_0\
        );

    \I__226\ : IoInMux
    port map (
            O => \N__2429\,
            I => \N__2426\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2426\,
            I => \N__2423\
        );

    \I__224\ : Span12Mux_s4_h
    port map (
            O => \N__2423\,
            I => \N__2420\
        );

    \I__223\ : Odrv12
    port map (
            O => \N__2420\,
            I => masterreset_c_i
        );

    \I__222\ : ClkMux
    port map (
            O => \N__2417\,
            I => \N__2414\
        );

    \I__221\ : GlobalMux
    port map (
            O => \N__2414\,
            I => \N__2411\
        );

    \I__220\ : gio2CtrlBuf
    port map (
            O => \N__2411\,
            I => \arse.un1_io_0_1_g\
        );

    \I__219\ : IoInMux
    port map (
            O => \N__2408\,
            I => \N__2405\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2405\,
            I => \N__2402\
        );

    \I__217\ : Span4Mux_s1_v
    port map (
            O => \N__2402\,
            I => \N__2399\
        );

    \I__216\ : Sp12to4
    port map (
            O => \N__2399\,
            I => \N__2396\
        );

    \I__215\ : Span12Mux_h
    port map (
            O => \N__2396\,
            I => \N__2393\
        );

    \I__214\ : Span12Mux_v
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__213\ : Span12Mux_v
    port map (
            O => \N__2390\,
            I => \N__2387\
        );

    \I__212\ : Odrv12
    port map (
            O => \N__2387\,
            I => \top_pll_nrtthrth.PLLOUTCORE\
        );

    \INVarse.divseven.dout_0C\ : INV
    port map (
            O => \INVarse.divseven.dout_0C_net\,
            I => \N__5906\
        );

    \INVarse.apuresetoutregC\ : INV
    port map (
            O => \INVarse.apuresetoutregC_net\,
            I => \N__5913\
        );

    \INVarse.apusynclatchedC\ : INV
    port map (
            O => \INVarse.apusynclatchedC_net\,
            I => \N__2417\
        );

    \INVarse.diveight.dout_0C\ : INV
    port map (
            O => \INVarse.diveight.dout_0C_net\,
            I => \N__5911\
        );

    \INVarse.doingsevenC\ : INV
    port map (
            O => \INVarse.doingsevenC_net\,
            I => \N__5903\
        );

    \INVarse.cpuclkresetC\ : INV
    port map (
            O => \INVarse.cpuclkresetC_net\,
            I => \N__5907\
        );

    \INVarse.cpuresetoutregC\ : INV
    port map (
            O => \INVarse.cpuresetoutregC_net\,
            I => \N__5902\
        );

    \INVarse.cpuresetcount_0C\ : INV
    port map (
            O => \INVarse.cpuresetcount_0C_net\,
            I => \N__5901\
        );

    \IN_MUX_bfv_21_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_12_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \arses.un2_counter_cry_8\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_27_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_27_8_0_\
        );

    \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2408\,
            GLOBALBUFFEROUTPUT => \PLLOUTCORE_g\
        );

    \arse.divseven.io_0_RNIIG08\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2456\,
            GLOBALBUFFEROUTPUT => \arse.un1_io_0_1_g\
        );

    \masterreset_ibuf_RNIKP26_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2429\,
            GLOBALBUFFEROUTPUT => masterreset_c_i_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \masterreset_ibuf_RNIKP26_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => masterreset_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.un3_counter_cry_1_c_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2493\,
            in2 => \N__2687\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \debouncedn.un3_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.un3_counter_cry_1_THRU_LUT4_0_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2601\,
            in2 => \_gnd_net_\,
            in3 => \N__2519\,
            lcout => \debouncedn.un3_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \debouncedn.un3_counter_cry_1\,
            carryout => \debouncedn.un3_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.un3_counter_cry_2_THRU_LUT4_0_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2654\,
            in2 => \_gnd_net_\,
            in3 => \N__2516\,
            lcout => \debouncedn.un3_counter_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \debouncedn.un3_counter_cry_2\,
            carryout => \debouncedn.un3_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_4_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__2476\,
            in1 => \N__4660\,
            in2 => \N__2627\,
            in3 => \N__2513\,
            lcout => \debouncedn.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.out_RNO_1_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2651\,
            in2 => \_gnd_net_\,
            in3 => \N__2600\,
            lcout => OPEN,
            ltout => \debouncedn.counter18_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.out_RNO_0_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2475\,
            in1 => \N__2684\,
            in2 => \N__2498\,
            in3 => \N__2494\,
            lcout => \debouncedn.out_cnv_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_1_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__2495\,
            in1 => \N__2685\,
            in2 => \N__4666\,
            in3 => \N__2626\,
            lcout => \debouncedn.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__4587\,
            in1 => \_gnd_net_\,
            in2 => \N__2720\,
            in3 => \N__2811\,
            lcout => \debounceconsolereset.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_RNIBTPA2_4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__2652\,
            in1 => \N__2602\,
            in2 => \N__2477\,
            in3 => \N__4586\,
            lcout => \debouncedn.counter_RNIBTPA2Z0Z_4\,
            ltout => \debouncedn.counter_RNIBTPA2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__4588\,
            in1 => \_gnd_net_\,
            in2 => \N__2690\,
            in3 => \N__2686\,
            lcout => \debouncedn.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_1_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__2810\,
            in1 => \N__2715\,
            in2 => \N__4663\,
            in3 => \N__2735\,
            lcout => \debounceconsolereset.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_RNO_1_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__2780\,
            in1 => \_gnd_net_\,
            in2 => \N__2842\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \debounceconsolereset.counter18_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_RNO_0_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2870\,
            in1 => \N__2714\,
            in2 => \N__2663\,
            in3 => \N__2734\,
            lcout => \debounceconsolereset.out_cnv_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_3_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__2621\,
            in1 => \N__2660\,
            in2 => \N__4638\,
            in3 => \N__2653\,
            lcout => \debouncedn.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.counter_2_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__2633\,
            in1 => \N__2603\,
            in2 => \N__4662\,
            in3 => \N__2622\,
            lcout => \debouncedn.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__2582\,
            in1 => \N__2561\,
            in2 => \N__6107\,
            in3 => \N__4637\,
            lcout => debouncedconsolereset,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \lcolreg_2_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4351\,
            in2 => \_gnd_net_\,
            in3 => \N__4488\,
            lcout => lcol3_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4780\,
            ce => \N__4682\,
            sr => \_gnd_net_\
        );

    \lcolreg_3_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4352\,
            in2 => \_gnd_net_\,
            in3 => \N__4489\,
            lcout => lcol4_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4780\,
            ce => \N__4682\,
            sr => \_gnd_net_\
        );

    \debounceup.un3_counter_cry_1_c_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2940\,
            in2 => \N__2993\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \debounceup.un3_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.un3_counter_cry_1_THRU_LUT4_0_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3028\,
            in2 => \_gnd_net_\,
            in3 => \N__2756\,
            lcout => \debounceup.un3_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceup.un3_counter_cry_1\,
            carryout => \debounceup.un3_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.un3_counter_cry_2_THRU_LUT4_0_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3049\,
            in2 => \_gnd_net_\,
            in3 => \N__2753\,
            lcout => \debounceup.un3_counter_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceup.un3_counter_cry_2\,
            carryout => \debounceup.un3_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_4_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__3011\,
            in1 => \N__4629\,
            in2 => \N__2969\,
            in3 => \N__2750\,
            lcout => \debounceup.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_3_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__2960\,
            in1 => \N__2747\,
            in2 => \N__4665\,
            in3 => \N__3050\,
            lcout => \debounceup.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_2_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__2741\,
            in1 => \N__3029\,
            in2 => \N__4664\,
            in3 => \N__2961\,
            lcout => \debounceup.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_1_c_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2733\,
            in2 => \N__2719\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \debounceconsolereset.un3_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2781\,
            in2 => \_gnd_net_\,
            in3 => \N__2696\,
            lcout => \debounceconsolereset.un3_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_1\,
            carryout => \debounceconsolereset.un3_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2843\,
            in3 => \N__2693\,
            lcout => \debounceconsolereset.un3_counter_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_2\,
            carryout => \debounceconsolereset.un3_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_4_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__2869\,
            in1 => \N__4618\,
            in2 => \N__2816\,
            in3 => \N__2873\,
            lcout => \debounceconsolereset.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_0_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__3559\,
            in1 => \N__3811\,
            in2 => \_gnd_net_\,
            in3 => \N__3397\,
            lcout => \clock_out_RNIR6ER_0\,
            ltout => \clock_out_RNIR6ER_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNINST81_4_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__2868\,
            in1 => \N__2837\,
            in2 => \N__2855\,
            in3 => \N__2782\,
            lcout => \debounceconsolereset.counter_RNINST81Z0Z_4\,
            ltout => \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_3_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4617\,
            in1 => \N__2852\,
            in2 => \N__2846\,
            in3 => \N__2841\,
            lcout => \debounceconsolereset.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_2_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__2783\,
            in1 => \N__2815\,
            in2 => \N__2792\,
            in3 => \N__4619\,
            lcout => \debounceconsolereset.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.un2_counter_cry_1_c_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3254\,
            in2 => \N__3116\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \arses.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_2_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3411\,
            in1 => \N__3134\,
            in2 => \_gnd_net_\,
            in3 => \N__2762\,
            lcout => \arses.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_1\,
            carryout => \arses.un2_counter_cry_2\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_3_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3405\,
            in1 => \N__3146\,
            in2 => \_gnd_net_\,
            in3 => \N__2759\,
            lcout => \arses.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_2\,
            carryout => \arses.un2_counter_cry_3\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_4_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3412\,
            in1 => \N__3266\,
            in2 => \_gnd_net_\,
            in3 => \N__2903\,
            lcout => \arses.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_3\,
            carryout => \arses.un2_counter_cry_4\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_5_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3406\,
            in1 => \N__3278\,
            in2 => \_gnd_net_\,
            in3 => \N__2900\,
            lcout => \arses.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_4\,
            carryout => \arses.un2_counter_cry_5\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_6_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3413\,
            in1 => \N__3305\,
            in2 => \_gnd_net_\,
            in3 => \N__2897\,
            lcout => \arses.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_5\,
            carryout => \arses.un2_counter_cry_6\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_7_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3407\,
            in1 => \N__3317\,
            in2 => \_gnd_net_\,
            in3 => \N__2894\,
            lcout => \arses.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_6\,
            carryout => \arses.un2_counter_cry_7\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_8_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3414\,
            in1 => \N__3292\,
            in2 => \_gnd_net_\,
            in3 => \N__2891\,
            lcout => \arses.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_7\,
            carryout => \arses.un2_counter_cry_8\,
            clk => \N__4768\,
            ce => 'H',
            sr => \N__4834\
        );

    \arses.counter_9_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3410\,
            in1 => \N__3200\,
            in2 => \_gnd_net_\,
            in3 => \N__2888\,
            lcout => \arses.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \arses.un2_counter_cry_9\,
            clk => \N__4774\,
            ce => 'H',
            sr => \N__4835\
        );

    \arses.counter_10_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3415\,
            in1 => \N__3215\,
            in2 => \_gnd_net_\,
            in3 => \N__2885\,
            lcout => \arses.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_9\,
            carryout => \arses.un2_counter_cry_10\,
            clk => \N__4774\,
            ce => 'H',
            sr => \N__4835\
        );

    \arses.counter_11_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3408\,
            in1 => \N__3227\,
            in2 => \_gnd_net_\,
            in3 => \N__2882\,
            lcout => \arses.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_10\,
            carryout => \arses.un2_counter_cry_11\,
            clk => \N__4774\,
            ce => 'H',
            sr => \N__4835\
        );

    \arses.counter_12_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3416\,
            in1 => \N__3161\,
            in2 => \_gnd_net_\,
            in3 => \N__2879\,
            lcout => \arses.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_11\,
            carryout => \arses.un2_counter_cry_12\,
            clk => \N__4774\,
            ce => 'H',
            sr => \N__4835\
        );

    \arses.counter_13_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3409\,
            in1 => \N__3176\,
            in2 => \_gnd_net_\,
            in3 => \N__2876\,
            lcout => \arses.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_12\,
            carryout => \arses.un2_counter_cry_13\,
            clk => \N__4774\,
            ce => 'H',
            sr => \N__4835\
        );

    \arses.counter_14_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3417\,
            in1 => \N__3188\,
            in2 => \_gnd_net_\,
            in3 => \N__3080\,
            lcout => \arses.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4774\,
            ce => 'H',
            sr => \N__4835\
        );

    \arses.counter_1_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3252\,
            in1 => \N__3112\,
            in2 => \_gnd_net_\,
            in3 => \N__3419\,
            lcout => \arses.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4779\,
            ce => 'H',
            sr => \N__4836\
        );

    \dig1.leds_1_i_3_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__5729\,
            in1 => \N__3485\,
            in2 => \N__5092\,
            in3 => \N__3086\,
            lcout => leds_1_i_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4761\,
            ce => \N__4680\,
            sr => \_gnd_net_\
        );

    \debounceup.counter_RNI45V02_4_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__3048\,
            in1 => \N__3009\,
            in2 => \N__4639\,
            in3 => \N__3027\,
            lcout => \debounceup.counter_RNI45V02Z0Z_4\,
            ltout => \debounceup.counter_RNI45V02Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_0_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4595\,
            in2 => \N__3053\,
            in3 => \N__2988\,
            lcout => \debounceup.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.out_RNO_1_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3047\,
            in2 => \_gnd_net_\,
            in3 => \N__3026\,
            lcout => OPEN,
            ltout => \debounceup.counter18_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.out_RNO_0_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3010\,
            in1 => \N__2984\,
            in2 => \N__2996\,
            in3 => \N__2941\,
            lcout => \debounceup.out_cnv_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.counter_1_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__2942\,
            in1 => \N__4633\,
            in2 => \N__2992\,
            in3 => \N__2965\,
            lcout => \debounceup.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_2_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000011"
        )
    port map (
            in0 => \N__3425\,
            in1 => \N__3443\,
            in2 => \N__5737\,
            in3 => \N__3431\,
            lcout => leds_1_i_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4770\,
            ce => \N__4681\,
            sr => \_gnd_net_\
        );

    \arses.counter_RNIA58_5_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3316\,
            in1 => \N__3304\,
            in2 => \N__3293\,
            in3 => \N__3277\,
            lcout => OPEN,
            ltout => \arses.un1_counterlto8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOKH_1_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3265\,
            in1 => \N__3253\,
            in2 => \N__3230\,
            in3 => \N__3122\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI04C4_9_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3226\,
            in1 => \N__3214\,
            in2 => \N__3203\,
            in3 => \N__3199\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOS0A_14_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__3187\,
            in1 => \N__3175\,
            in2 => \N__3164\,
            in3 => \N__3160\,
            lcout => \arses.counter8\,
            ltout => \arses.counter8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__3584\,
            in1 => \_gnd_net_\,
            in2 => \N__3149\,
            in3 => \N__3819\,
            lcout => slowclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI1L5_2_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3145\,
            in1 => \N__3133\,
            in2 => \_gnd_net_\,
            in3 => \N__3107\,
            lcout => \arses.un1_counterlto4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_0_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3111\,
            in2 => \_gnd_net_\,
            in3 => \N__3418\,
            lcout => \arses.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4782\,
            ce => 'H',
            sr => \N__4837\
        );

    \dig1.leds_cnst_3_1__m77_ns_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3677\,
            in1 => \N__3728\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \dig1.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m71_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001000000"
        )
    port map (
            in0 => \N__4201\,
            in1 => \N__5506\,
            in2 => \N__4490\,
            in3 => \N__4349\,
            lcout => \dig1.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.out_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__3479\,
            in1 => \N__3467\,
            in2 => \N__3509\,
            in3 => \N__4678\,
            lcout => debounceddn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m57_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111010010"
        )
    port map (
            in0 => \N__4334\,
            in1 => \N__5496\,
            in2 => \N__4216\,
            in3 => \N__4454\,
            lcout => OPEN,
            ltout => \dig1.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__3437\,
            in1 => \N__5728\,
            in2 => \N__3446\,
            in3 => \N__5087\,
            lcout => \dig1.leds_17_i_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m60_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110110100000"
        )
    port map (
            in0 => \N__4333\,
            in1 => \N__5495\,
            in2 => \N__4215\,
            in3 => \N__4453\,
            lcout => \dig1.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m68_bm_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111010010010"
        )
    port map (
            in0 => \N__4466\,
            in1 => \N__4212\,
            in2 => \N__5512\,
            in3 => \N__4115\,
            lcout => \dig1.m68_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m68_am_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010001000"
        )
    port map (
            in0 => \N__4322\,
            in1 => \N__5502\,
            in2 => \N__4217\,
            in3 => \N__4465\,
            lcout => \dig1.m68_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__3812\,
            in1 => \N__3583\,
            in2 => \_gnd_net_\,
            in3 => \N__3398\,
            lcout => \clock_out_RNIR6ER\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \lcolreg_1_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4330\,
            in2 => \_gnd_net_\,
            in3 => \N__4471\,
            lcout => lcol2_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4783\,
            ce => \N__4690\,
            sr => \_gnd_net_\
        );

    \delayConstant_0_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__3912\,
            in1 => \N__3874\,
            in2 => \_gnd_net_\,
            in3 => \N__5708\,
            lcout => \delayConstantZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4762\,
            ce => 'H',
            sr => \N__4839\
        );

    \olddn_RNIM5BH1_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3907\,
            in2 => \_gnd_net_\,
            in3 => \N__3868\,
            lcout => \olddn_RNIM5BHZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oldup_RNI8NJV_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__3585\,
            in1 => \N__3515\,
            in2 => \_gnd_net_\,
            in3 => \N__3690\,
            lcout => \delayConstant16_i\,
            ltout => \delayConstant16_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_0_c_RNO_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \N__5712\,
            in1 => \_gnd_net_\,
            in2 => \N__3518\,
            in3 => \N__3867\,
            lcout => \un1_delayConstant_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_3_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__3869\,
            in1 => \_gnd_net_\,
            in2 => \N__3914\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNIM5BH1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIEENH_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3491\,
            in2 => \_gnd_net_\,
            in3 => \N__3504\,
            lcout => \olddn_RNIEENHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oldup_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3691\,
            lcout => \oldupZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_0_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3911\,
            in2 => \_gnd_net_\,
            in3 => \N__3870\,
            lcout => \olddn_RNIM5BH1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \olddnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m77_am_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001110101011"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__4172\,
            in2 => \N__5493\,
            in3 => \N__4473\,
            lcout => \dig1.m77_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.out_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__3722\,
            in1 => \N__3692\,
            in2 => \N__3710\,
            in3 => \N__4679\,
            lcout => debouncedup,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m77_bm_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4472\,
            in1 => \N__4331\,
            in2 => \N__4197\,
            in3 => \N__5466\,
            lcout => \dig1.m77_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m35_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000001000"
        )
    port map (
            in0 => \N__4335\,
            in1 => \N__5385\,
            in2 => \N__4050\,
            in3 => \N__4474\,
            lcout => \dig1.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_1_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3830\,
            in1 => \N__4058\,
            in2 => \_gnd_net_\,
            in3 => \N__5779\,
            lcout => leds_1_i_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4781\,
            ce => \N__4694\,
            sr => \_gnd_net_\
        );

    \lcolreg_0_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4329\,
            in2 => \_gnd_net_\,
            in3 => \N__4470\,
            lcout => lcol1_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4781\,
            ce => \N__4694\,
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_3_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__4067\,
            in1 => \N__5780\,
            in2 => \N__5158\,
            in3 => \N__3632\,
            lcout => leds_1_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4781\,
            ce => \N__4694\,
            sr => \_gnd_net_\
        );

    \col_1_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__4311\,
            in1 => \N__4114\,
            in2 => \N__3824\,
            in3 => \N__3788\,
            lcout => \colZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m14_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100010101"
        )
    port map (
            in0 => \N__4047\,
            in1 => \N__4310\,
            in2 => \N__5417\,
            in3 => \N__4449\,
            lcout => OPEN,
            ltout => \dig1.N_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m17_ns_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3779\,
            in2 => \N__3833\,
            in3 => \N__5154\,
            lcout => \dig1.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \col_0_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__4450\,
            in1 => \N__3820\,
            in2 => \_gnd_net_\,
            in3 => \N__3787\,
            lcout => \colZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m16_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000010010"
        )
    port map (
            in0 => \N__4046\,
            in1 => \N__4309\,
            in2 => \N__5416\,
            in3 => \N__4448\,
            lcout => \dig1.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m32_am_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000001000"
        )
    port map (
            in0 => \N__4052\,
            in1 => \N__4464\,
            in2 => \N__4350\,
            in3 => \N__5405\,
            lcout => \dig1.m32_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m32_bm_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111010010010"
        )
    port map (
            in0 => \N__4463\,
            in1 => \N__4051\,
            in2 => \N__5418\,
            in3 => \N__4113\,
            lcout => \dig1.m32_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_2_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001010101"
        )
    port map (
            in0 => \N__4871\,
            in1 => \N__3773\,
            in2 => \N__3767\,
            in3 => \N__5785\,
            lcout => leds_1_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4786\,
            ce => \N__4689\,
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_1_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3904\,
            in2 => \_gnd_net_\,
            in3 => \N__3871\,
            lcout => \olddn_RNIM5BH1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_4_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3906\,
            in2 => \_gnd_net_\,
            in3 => \N__3873\,
            lcout => \olddn_RNIM5BH1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNIM5BH1_2_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3905\,
            in2 => \_gnd_net_\,
            in3 => \N__3872\,
            lcout => \olddn_RNIM5BH1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_0_c_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5697\,
            in2 => \N__3737\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_12_0_\,
            carryout => \un1_delayConstant_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_1_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3983\,
            in2 => \N__5494\,
            in3 => \N__3977\,
            lcout => \delayConstantZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_0\,
            carryout => \un1_delayConstant_cry_1\,
            clk => \N__4772\,
            ce => 'H',
            sr => \N__4840\
        );

    \un1_delayConstant_cry_1_0_c_RNIJGN92_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3974\,
            in2 => \N__4214\,
            in3 => \N__3968\,
            lcout => \un1_delayConstant_cry_1_0_c_RNIJGNZ0Z92\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_1\,
            carryout => \un1_delayConstant_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_3_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5058\,
            in2 => \N__3965\,
            in3 => \N__3956\,
            lcout => \delayConstantZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_2\,
            carryout => \un1_delayConstant_cry_3\,
            clk => \N__4772\,
            ce => 'H',
            sr => \N__4840\
        );

    \delayConstant_4_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5759\,
            in2 => \N__3953\,
            in3 => \N__3941\,
            lcout => \delayConstantZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_3\,
            carryout => \un1_delayConstant_cry_4\,
            clk => \N__4772\,
            ce => 'H',
            sr => \N__4840\
        );

    \delayConstant_5_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3938\,
            in2 => \N__5386\,
            in3 => \N__3932\,
            lcout => \delayConstantZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_4\,
            carryout => \un1_delayConstant_cry_5\,
            clk => \N__4772\,
            ce => 'H',
            sr => \N__4840\
        );

    \un1_delayConstant_cry_5_0_c_RNIR4GA2_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4036\,
            in2 => \N__3929\,
            in3 => \N__3917\,
            lcout => \un1_delayConstant_cry_5_0_c_RNIR4GAZ0Z2\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_5\,
            carryout => \un1_delayConstant_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_7_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__3913\,
            in1 => \N__3875\,
            in2 => \N__5153\,
            in3 => \N__3836\,
            lcout => \delayConstantZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4772\,
            ce => 'H',
            sr => \N__4840\
        );

    \delayConstant_6_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4864\,
            lcout => \delayConstantZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4778\,
            ce => 'H',
            sr => \N__4838\
        );

    \delayConstant_2_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4852\,
            lcout => \delayConstantZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4778\,
            ce => 'H',
            sr => \N__4838\
        );

    \dig1.leds_cnst_3_1__m41_bm_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4039\,
            in1 => \N__4312\,
            in2 => \N__5406\,
            in3 => \N__4451\,
            lcout => \dig1.m41_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m41_am_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010111001101"
        )
    port map (
            in0 => \N__4040\,
            in1 => \N__4313\,
            in2 => \N__5407\,
            in3 => \N__4452\,
            lcout => OPEN,
            ltout => \dig1.m41_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m41_ns_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4076\,
            in2 => \N__4070\,
            in3 => \N__5147\,
            lcout => \dig1.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m2_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__4305\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4443\,
            lcout => col_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m10_ns_1_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__4445\,
            in1 => \N__4048\,
            in2 => \N__5419\,
            in3 => \N__4306\,
            lcout => OPEN,
            ltout => \dig1.m10_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m10_ns_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__4049\,
            in1 => \N__4112\,
            in2 => \N__4061\,
            in3 => \N__5152\,
            lcout => \dig1.N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m52_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000110010000"
        )
    port map (
            in0 => \N__4444\,
            in1 => \N__4304\,
            in2 => \N__4208\,
            in3 => \N__5489\,
            lcout => \dig1.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m24_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001110001000"
        )
    port map (
            in0 => \N__4037\,
            in1 => \N__4307\,
            in2 => \N__5414\,
            in3 => \N__4446\,
            lcout => \dig1.N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m21_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110100110"
        )
    port map (
            in0 => \N__4038\,
            in1 => \N__4308\,
            in2 => \N__5415\,
            in3 => \N__4447\,
            lcout => OPEN,
            ltout => \dig1.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__4880\,
            in1 => \N__5784\,
            in2 => \N__4874\,
            in3 => \N__5151\,
            lcout => \dig1.leds_17_i_0_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_fast_6_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4865\,
            lcout => \delayConstant_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4773\,
            ce => 'H',
            sr => \N__4841\
        );

    \delayConstant_fast_2_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \delayConstant_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4773\,
            ce => 'H',
            sr => \N__4841\
        );

    \dig1.leds_1_i_1_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4496\,
            in1 => \N__4082\,
            in2 => \_gnd_net_\,
            in3 => \N__5733\,
            lcout => leds_1_i_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4785\,
            ce => \N__4661\,
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m50_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100000111"
        )
    port map (
            in0 => \N__4336\,
            in1 => \N__5508\,
            in2 => \N__4213\,
            in3 => \N__4476\,
            lcout => OPEN,
            ltout => \dig1.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m53_ns_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5082\,
            in2 => \N__4505\,
            in3 => \N__4502\,
            lcout => \dig1.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m47_ns_1_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__4475\,
            in1 => \N__4195\,
            in2 => \N__5513\,
            in3 => \N__4337\,
            lcout => OPEN,
            ltout => \dig1.m47_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m47_ns_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__5083\,
            in1 => \N__4196\,
            in2 => \N__4118\,
            in3 => \N__4111\,
            lcout => \dig1.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_23_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_4_LC_27_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__5279\,
            in1 => \N__5660\,
            in2 => \N__5639\,
            in3 => \N__5306\,
            lcout => \arse.g0_i_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_0_LC_27_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5662\,
            in2 => \N__6194\,
            in3 => \N__6190\,
            lcout => \arse.cpuresetcountZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_27_8_0_\,
            carryout => \arse.un1_cpuresetcount_1_cry_0\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_1_LC_27_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5282\,
            in2 => \_gnd_net_\,
            in3 => \N__4898\,
            lcout => \arse.cpuresetcountZ0Z_1\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_0\,
            carryout => \arse.un1_cpuresetcount_1_cry_1\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_2_LC_27_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5181\,
            in2 => \_gnd_net_\,
            in3 => \N__4895\,
            lcout => \arse.cpuresetcountZ0Z_2\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_1\,
            carryout => \arse.un1_cpuresetcount_1_cry_2\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_3_LC_27_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4997\,
            in2 => \_gnd_net_\,
            in3 => \N__4892\,
            lcout => \arse.cpuresetcountZ0Z_3\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_2\,
            carryout => \arse.un1_cpuresetcount_1_cry_3\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_4_LC_27_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5638\,
            in2 => \_gnd_net_\,
            in3 => \N__4889\,
            lcout => \arse.cpuresetcountZ0Z_4\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_3\,
            carryout => \arse.un1_cpuresetcount_1_cry_4\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_5_LC_27_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5309\,
            in2 => \_gnd_net_\,
            in3 => \N__4886\,
            lcout => \arse.cpuresetcountZ0Z_5\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_4\,
            carryout => \arse.un1_cpuresetcount_1_cry_5\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_6_LC_27_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5210\,
            in2 => \_gnd_net_\,
            in3 => \N__4883\,
            lcout => \arse.cpuresetcountZ0Z_6\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_5\,
            carryout => \arse.un1_cpuresetcount_1_cry_6\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetcount_7_LC_27_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5020\,
            in2 => \_gnd_net_\,
            in3 => \N__5516\,
            lcout => \arse.cpuresetcountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5548\
        );

    \arse.cpuresetoutreg_RNO_2_LC_27_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__5507\,
            in1 => \N__5281\,
            in2 => \N__5423\,
            in3 => \N__5307\,
            lcout => \arse.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_1_LC_28_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5016\,
            in1 => \N__4994\,
            in2 => \N__5212\,
            in3 => \N__5315\,
            lcout => \arse.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_RNIATKJ1_7_LC_28_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5015\,
            in1 => \N__5308\,
            in2 => \N__5211\,
            in3 => \N__5636\,
            lcout => \arse.doingseven3_6\,
            ltout => \arse.doingseven3_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.doingseven_RNO_0_LC_28_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4996\,
            in1 => \N__5258\,
            in2 => \N__5285\,
            in3 => \N__5183\,
            lcout => \arse.doingseven3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_RNIB4QP_0_LC_28_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5280\,
            in2 => \_gnd_net_\,
            in3 => \N__5661\,
            lcout => \arse.doingseven3_1\,
            ltout => \arse.doingseven3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuclkreset_RNO_0_LC_28_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__4995\,
            in1 => \N__5252\,
            in2 => \N__5246\,
            in3 => \N__5182\,
            lcout => \arse.doingseven4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_7_LC_28_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__5243\,
            in1 => \N__5228\,
            in2 => \N__5213\,
            in3 => \N__5180\,
            lcout => \arse.g0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_6_LC_28_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__5162\,
            in1 => \N__5093\,
            in2 => \N__5021\,
            in3 => \N__4993\,
            lcout => \arse.g0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_5_LC_28_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__5786\,
            in1 => \N__5738\,
            in2 => \N__5669\,
            in3 => \N__5637\,
            lcout => OPEN,
            ltout => \arse.g0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_3_LC_28_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5612\,
            in2 => \N__5606\,
            in3 => \N__5603\,
            lcout => OPEN,
            ltout => \arse.g0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_0_LC_28_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__5591\,
            in2 => \N__5585\,
            in3 => \N__6189\,
            lcout => OPEN,
            ltout => \arse.cpuresetoutreg_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_LC_28_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5582\,
            in3 => \N__5575\,
            lcout => \arse.cpuresetoutregZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuresetoutregC_net\,
            ce => 'H',
            sr => \N__5547\
        );

    \arse.cpuclkreset_LC_29_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__6178\,
            in1 => \N__6048\,
            in2 => \_gnd_net_\,
            in3 => \N__5561\,
            lcout => \arse.cpuclkresetZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuclkresetC_net\,
            ce => 'H',
            sr => \N__5549\
        );

    \arse.doingseven_LC_29_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__6179\,
            in1 => \N__5818\,
            in2 => \_gnd_net_\,
            in3 => \N__5555\,
            lcout => \arse.doingsevenZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.doingsevenC_net\,
            ce => 'H',
            sr => \N__5540\
        );

    \debounceconsolereset.out_RNI1B6C_LC_29_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => debouncedconsolereset_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_0_LC_30_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6065\,
            in2 => \_gnd_net_\,
            in3 => \N__6039\,
            lcout => \arse.diveight.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_2_LC_30_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010000000"
        )
    port map (
            in0 => \N__6041\,
            in1 => \N__6010\,
            in2 => \N__6073\,
            in3 => \N__5992\,
            lcout => \arse.diveight.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_1_LC_30_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__6009\,
            in1 => \N__6066\,
            in2 => \_gnd_net_\,
            in3 => \N__6040\,
            lcout => \arse.diveight.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.seven_LC_30_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011000100"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__6232\,
            in2 => \N__5819\,
            in3 => \N__6264\,
            lcout => \arse.divseven.sevenZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_0_LC_31_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6050\,
            in2 => \_gnd_net_\,
            in3 => \N__5991\,
            lcout => \arse.diveight.doutZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.diveight.dout_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.seven_RNO_0_LC_31_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5859\,
            in2 => \_gnd_net_\,
            in3 => \N__5952\,
            lcout => \arse.divseven.un1_counter_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_0_LC_31_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__5860\,
            in1 => \N__5953\,
            in2 => \N__6265\,
            in3 => \N__6230\,
            lcout => \arse.divseven.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_2_LC_31_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111111000000"
        )
    port map (
            in0 => \N__6229\,
            in1 => \N__6257\,
            in2 => \N__5960\,
            in3 => \N__5862\,
            lcout => \arse.divseven.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_1_LC_31_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010000111100"
        )
    port map (
            in0 => \N__5861\,
            in1 => \N__5954\,
            in2 => \N__6266\,
            in3 => \N__6231\,
            lcout => \arse.divseven.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_RNO_0_1_LC_31_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__6256\,
            in1 => \_gnd_net_\,
            in2 => \N__6233\,
            in3 => \_gnd_net_\,
            lcout => \arse.divseven.N_46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_RNO_0_LC_31_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5858\,
            in1 => \N__6255\,
            in2 => \N__5959\,
            in3 => \N__6225\,
            lcout => \arse.divseven.un1_dout_2_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.apusynclatched_LC_32_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__6153\,
            in1 => \N__6206\,
            in2 => \_gnd_net_\,
            in3 => \N__6132\,
            lcout => \arse.apusynclatchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.apusynclatchedC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.apuresetoutreg_LC_32_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6140\,
            lcout => \arse.apuresetoutregZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.apuresetoutregC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_1_LC_32_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__6074\,
            in1 => \N__6049\,
            in2 => \N__6017\,
            in3 => \N__5996\,
            lcout => \arse.diveight.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_1_LC_32_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011110011001100"
        )
    port map (
            in0 => \N__5927\,
            in1 => \N__5864\,
            in2 => \N__5969\,
            in3 => \N__5958\,
            lcout => \arse.divseven.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_0_LC_32_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \arse.divseven.doutZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.divseven.dout_0C_net\,
            ce => \N__5828\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
