// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Nov 8 2023 16:58:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top_pll" view "INTERFACE"

module top_pll (
    led6,
    led2,
    lcol1,
    RESET,
    led7,
    led3,
    lcol4,
    PLLOUTCORE,
    PACKAGEPIN,
    led8,
    led4,
    lcol3,
    led5,
    led1,
    lcol2,
    PLLOUTGLOBAL);

    output led6;
    output led2;
    output lcol1;
    input RESET;
    output led7;
    output led3;
    output lcol4;
    output PLLOUTCORE;
    input PACKAGEPIN;
    output led8;
    output led4;
    output lcol3;
    output led5;
    output led1;
    output lcol2;
    output PLLOUTGLOBAL;

    wire N__3086;
    wire N__3072;
    wire N__3071;
    wire N__3070;
    wire N__3063;
    wire N__3062;
    wire N__3061;
    wire N__3054;
    wire N__3053;
    wire N__3052;
    wire N__3045;
    wire N__3044;
    wire N__3043;
    wire N__3036;
    wire N__3035;
    wire N__3034;
    wire N__3027;
    wire N__3026;
    wire N__3025;
    wire N__3018;
    wire N__3017;
    wire N__3016;
    wire N__3009;
    wire N__3008;
    wire N__3007;
    wire N__3000;
    wire N__2999;
    wire N__2998;
    wire N__2991;
    wire N__2990;
    wire N__2989;
    wire N__2982;
    wire N__2981;
    wire N__2980;
    wire N__2973;
    wire N__2972;
    wire N__2971;
    wire N__2964;
    wire N__2963;
    wire N__2962;
    wire N__2955;
    wire N__2954;
    wire N__2953;
    wire N__2946;
    wire N__2945;
    wire N__2944;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2908;
    wire N__2907;
    wire N__2906;
    wire N__2905;
    wire N__2902;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2860;
    wire N__2857;
    wire N__2856;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2824;
    wire N__2821;
    wire N__2820;
    wire N__2819;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2804;
    wire N__2801;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2779;
    wire N__2778;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2770;
    wire N__2769;
    wire N__2766;
    wire N__2765;
    wire N__2762;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2737;
    wire N__2726;
    wire N__2723;
    wire N__2722;
    wire N__2719;
    wire N__2718;
    wire N__2717;
    wire N__2716;
    wire N__2715;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2703;
    wire N__2700;
    wire N__2695;
    wire N__2684;
    wire N__2683;
    wire N__2682;
    wire N__2681;
    wire N__2680;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2665;
    wire N__2662;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2644;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2621;
    wire N__2620;
    wire N__2619;
    wire N__2618;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2606;
    wire N__2603;
    wire N__2594;
    wire N__2591;
    wire N__2590;
    wire N__2589;
    wire N__2588;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2576;
    wire N__2573;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2548;
    wire N__2545;
    wire N__2542;
    wire N__2541;
    wire N__2540;
    wire N__2535;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2505;
    wire N__2500;
    wire N__2499;
    wire N__2494;
    wire N__2491;
    wire N__2488;
    wire N__2485;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2467;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2450;
    wire N__2449;
    wire N__2448;
    wire N__2447;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2435;
    wire N__2432;
    wire N__2423;
    wire N__2422;
    wire N__2421;
    wire N__2420;
    wire N__2417;
    wire N__2416;
    wire N__2413;
    wire N__2410;
    wire N__2407;
    wire N__2404;
    wire N__2401;
    wire N__2398;
    wire N__2387;
    wire N__2386;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2376;
    wire N__2369;
    wire N__2368;
    wire N__2367;
    wire N__2366;
    wire N__2365;
    wire N__2362;
    wire N__2357;
    wire N__2352;
    wire N__2345;
    wire N__2344;
    wire N__2343;
    wire N__2342;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2327;
    wire N__2318;
    wire N__2317;
    wire N__2316;
    wire N__2315;
    wire N__2314;
    wire N__2311;
    wire N__2308;
    wire N__2303;
    wire N__2298;
    wire N__2291;
    wire N__2290;
    wire N__2287;
    wire N__2286;
    wire N__2285;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2271;
    wire N__2264;
    wire N__2261;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2251;
    wire N__2246;
    wire N__2245;
    wire N__2242;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2219;
    wire N__2216;
    wire N__2215;
    wire N__2212;
    wire N__2209;
    wire N__2206;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2187;
    wire N__2184;
    wire N__2181;
    wire N__2174;
    wire N__2173;
    wire N__2172;
    wire N__2169;
    wire N__2166;
    wire N__2163;
    wire N__2156;
    wire N__2155;
    wire N__2154;
    wire N__2153;
    wire N__2152;
    wire N__2149;
    wire N__2144;
    wire N__2139;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2123;
    wire N__2122;
    wire N__2119;
    wire N__2118;
    wire N__2117;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2105;
    wire N__2102;
    wire N__2093;
    wire N__2090;
    wire N__2087;
    wire N__2086;
    wire N__2085;
    wire N__2084;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2069;
    wire N__2066;
    wire N__2057;
    wire N__2054;
    wire N__2051;
    wire N__2048;
    wire N__2045;
    wire N__2042;
    wire N__2039;
    wire N__2038;
    wire N__2037;
    wire N__2036;
    wire N__2035;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2017;
    wire N__2016;
    wire N__2013;
    wire N__2010;
    wire N__2007;
    wire N__2000;
    wire N__1999;
    wire N__1996;
    wire N__1993;
    wire N__1988;
    wire N__1987;
    wire N__1984;
    wire N__1981;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1967;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1952;
    wire N__1949;
    wire N__1948;
    wire N__1945;
    wire N__1942;
    wire N__1941;
    wire N__1938;
    wire N__1935;
    wire N__1932;
    wire N__1925;
    wire N__1922;
    wire N__1919;
    wire N__1918;
    wire N__1915;
    wire N__1912;
    wire N__1907;
    wire N__1904;
    wire N__1903;
    wire N__1900;
    wire N__1897;
    wire N__1896;
    wire N__1891;
    wire N__1888;
    wire N__1885;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1871;
    wire N__1868;
    wire N__1867;
    wire N__1866;
    wire N__1865;
    wire N__1864;
    wire N__1863;
    wire N__1862;
    wire N__1861;
    wire N__1860;
    wire N__1857;
    wire N__1838;
    wire N__1835;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1817;
    wire N__1814;
    wire N__1811;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1796;
    wire N__1793;
    wire N__1790;
    wire N__1787;
    wire N__1784;
    wire N__1781;
    wire N__1778;
    wire N__1775;
    wire N__1772;
    wire N__1769;
    wire N__1766;
    wire N__1763;
    wire N__1760;
    wire N__1757;
    wire N__1754;
    wire N__1751;
    wire N__1748;
    wire N__1745;
    wire N__1742;
    wire N__1739;
    wire N__1736;
    wire N__1733;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1711;
    wire N__1710;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1695;
    wire N__1692;
    wire N__1689;
    wire N__1682;
    wire N__1681;
    wire N__1678;
    wire N__1677;
    wire N__1674;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1656;
    wire N__1653;
    wire N__1646;
    wire N__1645;
    wire N__1644;
    wire N__1643;
    wire N__1642;
    wire N__1639;
    wire N__1636;
    wire N__1629;
    wire N__1626;
    wire N__1623;
    wire N__1616;
    wire N__1613;
    wire N__1610;
    wire N__1607;
    wire N__1604;
    wire N__1603;
    wire N__1602;
    wire N__1601;
    wire N__1600;
    wire N__1599;
    wire N__1598;
    wire N__1597;
    wire N__1580;
    wire N__1579;
    wire N__1578;
    wire N__1577;
    wire N__1574;
    wire N__1571;
    wire N__1568;
    wire N__1565;
    wire N__1556;
    wire N__1555;
    wire N__1554;
    wire N__1553;
    wire N__1550;
    wire N__1547;
    wire N__1544;
    wire N__1543;
    wire N__1542;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1520;
    wire N__1519;
    wire N__1516;
    wire N__1515;
    wire N__1514;
    wire N__1513;
    wire N__1506;
    wire N__1503;
    wire N__1500;
    wire N__1493;
    wire N__1492;
    wire N__1491;
    wire N__1490;
    wire N__1489;
    wire N__1482;
    wire N__1479;
    wire N__1476;
    wire N__1469;
    wire N__1466;
    wire N__1463;
    wire N__1460;
    wire N__1459;
    wire N__1456;
    wire N__1453;
    wire N__1448;
    wire N__1445;
    wire N__1442;
    wire N__1439;
    wire N__1436;
    wire N__1433;
    wire N__1430;
    wire N__1427;
    wire N__1424;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1414;
    wire N__1411;
    wire N__1408;
    wire N__1403;
    wire N__1400;
    wire N__1397;
    wire N__1394;
    wire N__1391;
    wire N__1388;
    wire N__1385;
    wire N__1384;
    wire N__1381;
    wire N__1378;
    wire N__1373;
    wire N__1372;
    wire N__1369;
    wire N__1366;
    wire N__1365;
    wire N__1360;
    wire N__1357;
    wire N__1352;
    wire N__1349;
    wire N__1348;
    wire N__1345;
    wire N__1342;
    wire N__1337;
    wire N__1334;
    wire N__1331;
    wire N__1328;
    wire N__1325;
    wire N__1322;
    wire N__1319;
    wire N__1316;
    wire N__1315;
    wire N__1312;
    wire N__1309;
    wire N__1306;
    wire N__1303;
    wire N__1298;
    wire N__1295;
    wire N__1292;
    wire N__1289;
    wire N__1286;
    wire N__1283;
    wire N__1280;
    wire N__1277;
    wire N__1274;
    wire N__1271;
    wire N__1268;
    wire N__1265;
    wire N__1262;
    wire N__1259;
    wire VCCG0;
    wire RESET_c;
    wire PLLOUTCORE_c;
    wire GNDG0;
    wire GB_BUFFER_PLLOUTGLOBAL_0_THRU_CO;
    wire \II_2.outputsZ0Z_1 ;
    wire \II_2.outputsZ0Z_0 ;
    wire \II_1.g3_3_cascade_ ;
    wire \II_1.counter_RNIIPRU2Z0Z_11_cascade_ ;
    wire \II_1.g0_1_a4_0_0 ;
    wire II_1_un2_clock_outlt27_0_i;
    wire \II_3.outputsZ0Z_0 ;
    wire \II_3.o2_cascade_ ;
    wire \II_2.un1_counter23_1_5 ;
    wire \II_2.counterZ0Z_2 ;
    wire \II_2.counterZ0Z_0 ;
    wire \II_2.counterZ0Z_1 ;
    wire \II_2.un1_counter19_1_0 ;
    wire counter_RNI6D8K_6_cascade_;
    wire counter_RNI6D8K_6;
    wire \II_1.clock_out_RNOZ0Z_5_cascade_ ;
    wire \II_1.counter_RNIK1FB1Z0Z_13 ;
    wire \II_1.counter_RNIJLJ01_0Z0Z_17 ;
    wire \II_1.un1_counterlt12_2 ;
    wire \II_3.N_14 ;
    wire \II_3.G_30_0_o3_0_1_cascade_ ;
    wire \II_1.counter_RNI1TC9Z0Z_8 ;
    wire \II_3.N_16 ;
    wire \II_3.G_30_0_a3_1 ;
    wire \II_3.outputs_RNO_0Z0Z_0 ;
    wire \II_3.counterZ0Z_1 ;
    wire \II_3.counterZ0Z_2 ;
    wire \II_3.counterZ0Z_0 ;
    wire \II_3.o2_0_cascade_ ;
    wire \II_3.N_12 ;
    wire II_2_G_3_out;
    wire \II_3.G_30_0_o3_0 ;
    wire \II_1.counter_RNIM7JB1Z0Z_22_cascade_ ;
    wire \II_1.counter_RNI64GM1Z0Z_26 ;
    wire bfn_15_29_0_;
    wire \II_1.counter_1_cry_1 ;
    wire \II_1.counter_1_cry_2 ;
    wire \II_1.counter_1_cry_3 ;
    wire \II_1.counter_1_cry_4 ;
    wire \II_1.counter_1_cry_5 ;
    wire \II_1.counter_1_cry_6 ;
    wire \II_1.counter_1_cry_7 ;
    wire \II_1.counter_1_cry_8 ;
    wire bfn_15_30_0_;
    wire \II_1.counter_1_cry_9 ;
    wire \II_1.counter_1_cry_10 ;
    wire \II_1.counter_1_cry_11 ;
    wire \II_1.counter_1_cry_12 ;
    wire \II_1.counter_1_cry_13 ;
    wire \II_1.counter_1_cry_14 ;
    wire \II_1.counter_1_cry_15 ;
    wire \II_1.counter_1_cry_16 ;
    wire bfn_15_31_0_;
    wire \II_1.counter_1_cry_17 ;
    wire \II_1.counter_1_cry_18 ;
    wire \II_1.counter_1_cry_19 ;
    wire \II_1.counter_1_cry_20 ;
    wire \II_1.counter_1_cry_21 ;
    wire \II_1.counter_1_cry_22 ;
    wire \II_1.counter_1_cry_23 ;
    wire \II_1.counter_1_cry_24 ;
    wire bfn_15_32_0_;
    wire \II_1.counter_1_cry_25 ;
    wire \II_1.counter_1_cry_26 ;
    wire \II_1.un1_counter_0_g ;
    wire \II_1.counterZ0Z_6 ;
    wire \II_1.counterZ0Z_2 ;
    wire \II_1.counterZ0Z_3 ;
    wire \II_1.un2_clock_outlto19_1_cascade_ ;
    wire \II_1.un2_clock_outlto19_1 ;
    wire \II_1.clock_out_RNOZ0Z_3 ;
    wire \II_1.un2_clock_outlto23_0_0_d_1_cascade_ ;
    wire counter_RNIG1JB1_20;
    wire \II_1.un2_clock_outlto23_0_0_d_cascade_ ;
    wire led8_c;
    wire PLLOUTGLOBAL_0;
    wire \II_3.outputs_RNO_10Z0Z_0_cascade_ ;
    wire \II_3.G_30_0_a3_2_3 ;
    wire \II_1.counterZ0Z_10 ;
    wire II_1_counter_9;
    wire II_1_counter_11;
    wire \II_1.counterZ0Z_7 ;
    wire II_1_counter_16;
    wire II_1_counter_15;
    wire II_1_counter_17;
    wire II_1_counter_14;
    wire \II_1.counterZ0Z_4 ;
    wire \II_1.counterZ0Z_1 ;
    wire \II_1.counterZ0Z_5 ;
    wire \II_1.counterZ0Z_0 ;
    wire \II_1.counterZ0Z_21 ;
    wire II_1_counter_22;
    wire \II_1.un2_clock_outlto23_0_0_c ;
    wire II_1_counter_13;
    wire \II_1.counter_RNIQ7FB1Z0Z_14 ;
    wire II_1_counter_8;
    wire \II_1.counter_RNI6VAM1Z0Z_13_cascade_ ;
    wire \II_1.counter_RNIJ54VZ0Z_7 ;
    wire \II_1.counter_RNIA1PIZ0Z_1 ;
    wire \II_1.counter_RNIJS2EZ0Z_2 ;
    wire II_1_counter_12;
    wire \II_1.counter_RNI49153Z0Z_8 ;
    wire II_1_counter_27;
    wire \II_1.counter_RNICTOG4Z0Z_12_cascade_ ;
    wire \II_1.un1_counter_0 ;
    wire II_1_counter_26;
    wire \II_1.un1_counterlto22_0 ;
    wire \II_1.un1_counterlto24_0_0 ;
    wire II_1_counter_25;
    wire II_1_counter_24;
    wire II_1_counter_23;
    wire \II_1.un1_counterlto25 ;
    wire \II_1.counterZ0Z_20 ;
    wire II_1_counter_19;
    wire \II_1.un1_counterlto25_cascade_ ;
    wire II_1_counter_18;
    wire \II_1.counter_RNINVA12Z0Z_20 ;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam top_pll_inst_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam top_pll_inst_pll.TEST_MODE=1'b0;
    defparam top_pll_inst_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam top_pll_inst_pll.PLLOUT_SELECT="GENCLK";
    defparam top_pll_inst_pll.FILTER_RANGE=3'b001;
    defparam top_pll_inst_pll.FEEDBACK_PATH="SIMPLE";
    defparam top_pll_inst_pll.FDA_RELATIVE=4'b0000;
    defparam top_pll_inst_pll.FDA_FEEDBACK=4'b0000;
    defparam top_pll_inst_pll.ENABLE_ICEGATE=1'b0;
    defparam top_pll_inst_pll.DIVR=4'b0000;
    defparam top_pll_inst_pll.DIVQ=3'b010;
    defparam top_pll_inst_pll.DIVF=7'b0111000;
    defparam top_pll_inst_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 top_pll_inst_pll (
            .PLLOUTGLOBAL(PLLOUTGLOBAL_0),
            .SDI(),
            .BYPASS(GNDG0),
            .RESETB(N__1298),
            .PLLOUTCORE(PLLOUTCORE_c),
            .LOCK(),
            .SDO(),
            .SCLK(),
            .LATCHINPUTVALUE(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__3086));
    IO_PAD top_pll_inst_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__3086),
            .PACKAGEPIN(PACKAGEPIN));
    defparam \II_3.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \II_3.io_0_iopad .PULLUP=1'b0;
    IO_PAD \II_3.io_0_iopad  (
            .OE(N__3072),
            .DIN(N__3071),
            .DOUT(N__3070),
            .PACKAGEPIN(led6));
    defparam \II_3.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \II_3.io_0_preio  (
            .PADOEN(N__3072),
            .PADOUT(N__3071),
            .PADIN(N__3070),
            .CLOCKENABLE(),
            .DOUT1(N__1372),
            .OUTPUTENABLE(N__2541),
            .DIN0(),
            .DOUT0(N__1373),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1903));
    IO_PAD lcol1_obuf_iopad (
            .OE(N__3063),
            .DIN(N__3062),
            .DOUT(N__3061),
            .PACKAGEPIN(lcol1));
    defparam lcol1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol1_obuf_preio (
            .PADOEN(N__3063),
            .PADOUT(N__3062),
            .PADIN(N__3061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol3_obuf_iopad (
            .OE(N__3054),
            .DIN(N__3053),
            .DOUT(N__3052),
            .PACKAGEPIN(lcol3));
    defparam lcol3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol3_obuf_preio (
            .PADOEN(N__3054),
            .PADOUT(N__3053),
            .PADIN(N__3052),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2534),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led1_obuft_iopad (
            .OE(N__3045),
            .DIN(N__3044),
            .DOUT(N__3043),
            .PACKAGEPIN(led1));
    defparam led1_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led1_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led1_obuft_preio (
            .PADOEN(N__3045),
            .PADOUT(N__3044),
            .PADIN(N__3043),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PLLOUTGLOBAL_obuf_iopad (
            .OE(N__3036),
            .DIN(N__3035),
            .DOUT(N__3034),
            .PACKAGEPIN(PLLOUTGLOBAL));
    defparam PLLOUTGLOBAL_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PLLOUTGLOBAL_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PLLOUTGLOBAL_obuf_preio (
            .PADOEN(N__3036),
            .PADOUT(N__3035),
            .PADIN(N__3034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1337),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led2_obuft_iopad (
            .OE(N__3027),
            .DIN(N__3026),
            .DOUT(N__3025),
            .PACKAGEPIN(led2));
    defparam led2_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led2_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led2_obuft_preio (
            .PADOEN(N__3027),
            .PADOUT(N__3026),
            .PADIN(N__3025),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol4_obuf_iopad (
            .OE(N__3018),
            .DIN(N__3017),
            .DOUT(N__3016),
            .PACKAGEPIN(lcol4));
    defparam lcol4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol4_obuf_preio (
            .PADOEN(N__3018),
            .PADOUT(N__3017),
            .PADIN(N__3016),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2548),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led4_obuft_iopad (
            .OE(N__3009),
            .DIN(N__3008),
            .DOUT(N__3007),
            .PACKAGEPIN(led4));
    defparam led4_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led4_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led4_obuft_preio (
            .PADOEN(N__3009),
            .PADOUT(N__3008),
            .PADIN(N__3007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PLLOUTCORE_obuf_iopad (
            .OE(N__3000),
            .DIN(N__2999),
            .DOUT(N__2998),
            .PACKAGEPIN(PLLOUTCORE));
    defparam PLLOUTCORE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PLLOUTCORE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PLLOUTCORE_obuf_preio (
            .PADOEN(N__3000),
            .PADOUT(N__2999),
            .PADIN(N__2998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1280),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol2_obuf_iopad (
            .OE(N__2991),
            .DIN(N__2990),
            .DOUT(N__2989),
            .PACKAGEPIN(lcol2));
    defparam lcol2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol2_obuf_preio (
            .PADOEN(N__2991),
            .PADOUT(N__2990),
            .PADIN(N__2989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2499),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \II_2.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \II_2.io_0_iopad .PULLUP=1'b0;
    IO_PAD \II_2.io_0_iopad  (
            .OE(N__2982),
            .DIN(N__2981),
            .DOUT(N__2980),
            .PACKAGEPIN(led7));
    defparam \II_2.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \II_2.io_0_preio  (
            .PADOEN(N__2982),
            .PADOUT(N__2981),
            .PADIN(N__2980),
            .CLOCKENABLE(),
            .DOUT1(N__1325),
            .OUTPUTENABLE(N__2558),
            .DIN0(),
            .DOUT0(N__1427),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__1918));
    IO_PAD led8_obuf_iopad (
            .OE(N__2973),
            .DIN(N__2972),
            .DOUT(N__2971),
            .PACKAGEPIN(led8));
    defparam led8_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led8_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led8_obuf_preio (
            .PADOEN(N__2973),
            .PADOUT(N__2972),
            .PADIN(N__2971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1922),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led3_obuft_iopad (
            .OE(N__2964),
            .DIN(N__2963),
            .DOUT(N__2962),
            .PACKAGEPIN(led3));
    defparam led3_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led3_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led3_obuft_preio (
            .PADOEN(N__2964),
            .PADOUT(N__2963),
            .PADIN(N__2962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led5_obuft_iopad (
            .OE(N__2955),
            .DIN(N__2954),
            .DOUT(N__2953),
            .PACKAGEPIN(led5));
    defparam led5_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led5_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led5_obuft_preio (
            .PADOEN(N__2955),
            .PADOUT(N__2954),
            .PADIN(N__2953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESET_ibuf_iopad (
            .OE(N__2946),
            .DIN(N__2945),
            .DOUT(N__2944),
            .PACKAGEPIN(RESET));
    defparam RESET_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESET_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESET_ibuf_preio (
            .PADOEN(N__2946),
            .PADOUT(N__2945),
            .PADIN(N__2944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESET_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__665 (
            .O(N__2927),
            .I(N__2924));
    LocalMux I__664 (
            .O(N__2924),
            .I(\II_1.counter_RNIA1PIZ0Z_1 ));
    InMux I__663 (
            .O(N__2921),
            .I(N__2918));
    LocalMux I__662 (
            .O(N__2918),
            .I(N__2915));
    Odrv12 I__661 (
            .O(N__2915),
            .I(\II_1.counter_RNIJS2EZ0Z_2 ));
    CascadeMux I__660 (
            .O(N__2912),
            .I(N__2909));
    InMux I__659 (
            .O(N__2909),
            .I(N__2902));
    CascadeMux I__658 (
            .O(N__2908),
            .I(N__2898));
    InMux I__657 (
            .O(N__2907),
            .I(N__2895));
    InMux I__656 (
            .O(N__2906),
            .I(N__2892));
    InMux I__655 (
            .O(N__2905),
            .I(N__2889));
    LocalMux I__654 (
            .O(N__2902),
            .I(N__2886));
    InMux I__653 (
            .O(N__2901),
            .I(N__2883));
    InMux I__652 (
            .O(N__2898),
            .I(N__2880));
    LocalMux I__651 (
            .O(N__2895),
            .I(II_1_counter_12));
    LocalMux I__650 (
            .O(N__2892),
            .I(II_1_counter_12));
    LocalMux I__649 (
            .O(N__2889),
            .I(II_1_counter_12));
    Odrv4 I__648 (
            .O(N__2886),
            .I(II_1_counter_12));
    LocalMux I__647 (
            .O(N__2883),
            .I(II_1_counter_12));
    LocalMux I__646 (
            .O(N__2880),
            .I(II_1_counter_12));
    InMux I__645 (
            .O(N__2867),
            .I(N__2864));
    LocalMux I__644 (
            .O(N__2864),
            .I(\II_1.counter_RNI49153Z0Z_8 ));
    InMux I__643 (
            .O(N__2861),
            .I(N__2857));
    InMux I__642 (
            .O(N__2860),
            .I(N__2852));
    LocalMux I__641 (
            .O(N__2857),
            .I(N__2849));
    InMux I__640 (
            .O(N__2856),
            .I(N__2846));
    InMux I__639 (
            .O(N__2855),
            .I(N__2843));
    LocalMux I__638 (
            .O(N__2852),
            .I(II_1_counter_27));
    Odrv4 I__637 (
            .O(N__2849),
            .I(II_1_counter_27));
    LocalMux I__636 (
            .O(N__2846),
            .I(II_1_counter_27));
    LocalMux I__635 (
            .O(N__2843),
            .I(II_1_counter_27));
    CascadeMux I__634 (
            .O(N__2834),
            .I(\II_1.counter_RNICTOG4Z0Z_12_cascade_ ));
    IoInMux I__633 (
            .O(N__2831),
            .I(N__2828));
    LocalMux I__632 (
            .O(N__2828),
            .I(\II_1.un1_counter_0 ));
    InMux I__631 (
            .O(N__2825),
            .I(N__2821));
    CascadeMux I__630 (
            .O(N__2824),
            .I(N__2815));
    LocalMux I__629 (
            .O(N__2821),
            .I(N__2812));
    InMux I__628 (
            .O(N__2820),
            .I(N__2809));
    InMux I__627 (
            .O(N__2819),
            .I(N__2804));
    InMux I__626 (
            .O(N__2818),
            .I(N__2804));
    InMux I__625 (
            .O(N__2815),
            .I(N__2801));
    Odrv4 I__624 (
            .O(N__2812),
            .I(II_1_counter_26));
    LocalMux I__623 (
            .O(N__2809),
            .I(II_1_counter_26));
    LocalMux I__622 (
            .O(N__2804),
            .I(II_1_counter_26));
    LocalMux I__621 (
            .O(N__2801),
            .I(II_1_counter_26));
    InMux I__620 (
            .O(N__2792),
            .I(N__2789));
    LocalMux I__619 (
            .O(N__2789),
            .I(\II_1.un1_counterlto22_0 ));
    InMux I__618 (
            .O(N__2786),
            .I(N__2783));
    LocalMux I__617 (
            .O(N__2783),
            .I(\II_1.un1_counterlto24_0_0 ));
    InMux I__616 (
            .O(N__2780),
            .I(N__2774));
    InMux I__615 (
            .O(N__2779),
            .I(N__2771));
    InMux I__614 (
            .O(N__2778),
            .I(N__2766));
    CascadeMux I__613 (
            .O(N__2777),
            .I(N__2762));
    LocalMux I__612 (
            .O(N__2774),
            .I(N__2757));
    LocalMux I__611 (
            .O(N__2771),
            .I(N__2757));
    InMux I__610 (
            .O(N__2770),
            .I(N__2754));
    InMux I__609 (
            .O(N__2769),
            .I(N__2751));
    LocalMux I__608 (
            .O(N__2766),
            .I(N__2748));
    InMux I__607 (
            .O(N__2765),
            .I(N__2745));
    InMux I__606 (
            .O(N__2762),
            .I(N__2742));
    Span4Mux_v I__605 (
            .O(N__2757),
            .I(N__2737));
    LocalMux I__604 (
            .O(N__2754),
            .I(N__2737));
    LocalMux I__603 (
            .O(N__2751),
            .I(II_1_counter_25));
    Odrv4 I__602 (
            .O(N__2748),
            .I(II_1_counter_25));
    LocalMux I__601 (
            .O(N__2745),
            .I(II_1_counter_25));
    LocalMux I__600 (
            .O(N__2742),
            .I(II_1_counter_25));
    Odrv4 I__599 (
            .O(N__2737),
            .I(II_1_counter_25));
    CascadeMux I__598 (
            .O(N__2726),
            .I(N__2723));
    InMux I__597 (
            .O(N__2723),
            .I(N__2719));
    InMux I__596 (
            .O(N__2722),
            .I(N__2711));
    LocalMux I__595 (
            .O(N__2719),
            .I(N__2708));
    InMux I__594 (
            .O(N__2718),
            .I(N__2703));
    InMux I__593 (
            .O(N__2717),
            .I(N__2703));
    InMux I__592 (
            .O(N__2716),
            .I(N__2700));
    InMux I__591 (
            .O(N__2715),
            .I(N__2695));
    InMux I__590 (
            .O(N__2714),
            .I(N__2695));
    LocalMux I__589 (
            .O(N__2711),
            .I(II_1_counter_24));
    Odrv4 I__588 (
            .O(N__2708),
            .I(II_1_counter_24));
    LocalMux I__587 (
            .O(N__2703),
            .I(II_1_counter_24));
    LocalMux I__586 (
            .O(N__2700),
            .I(II_1_counter_24));
    LocalMux I__585 (
            .O(N__2695),
            .I(II_1_counter_24));
    InMux I__584 (
            .O(N__2684),
            .I(N__2676));
    InMux I__583 (
            .O(N__2683),
            .I(N__2673));
    InMux I__582 (
            .O(N__2682),
            .I(N__2670));
    InMux I__581 (
            .O(N__2681),
            .I(N__2665));
    InMux I__580 (
            .O(N__2680),
            .I(N__2665));
    InMux I__579 (
            .O(N__2679),
            .I(N__2662));
    LocalMux I__578 (
            .O(N__2676),
            .I(II_1_counter_23));
    LocalMux I__577 (
            .O(N__2673),
            .I(II_1_counter_23));
    LocalMux I__576 (
            .O(N__2670),
            .I(II_1_counter_23));
    LocalMux I__575 (
            .O(N__2665),
            .I(II_1_counter_23));
    LocalMux I__574 (
            .O(N__2662),
            .I(II_1_counter_23));
    InMux I__573 (
            .O(N__2651),
            .I(N__2648));
    LocalMux I__572 (
            .O(N__2648),
            .I(\II_1.un1_counterlto25 ));
    CascadeMux I__571 (
            .O(N__2645),
            .I(N__2640));
    InMux I__570 (
            .O(N__2644),
            .I(N__2637));
    InMux I__569 (
            .O(N__2643),
            .I(N__2634));
    InMux I__568 (
            .O(N__2640),
            .I(N__2631));
    LocalMux I__567 (
            .O(N__2637),
            .I(N__2628));
    LocalMux I__566 (
            .O(N__2634),
            .I(\II_1.counterZ0Z_20 ));
    LocalMux I__565 (
            .O(N__2631),
            .I(\II_1.counterZ0Z_20 ));
    Odrv4 I__564 (
            .O(N__2628),
            .I(\II_1.counterZ0Z_20 ));
    InMux I__563 (
            .O(N__2621),
            .I(N__2614));
    InMux I__562 (
            .O(N__2620),
            .I(N__2611));
    InMux I__561 (
            .O(N__2619),
            .I(N__2606));
    InMux I__560 (
            .O(N__2618),
            .I(N__2606));
    InMux I__559 (
            .O(N__2617),
            .I(N__2603));
    LocalMux I__558 (
            .O(N__2614),
            .I(II_1_counter_19));
    LocalMux I__557 (
            .O(N__2611),
            .I(II_1_counter_19));
    LocalMux I__556 (
            .O(N__2606),
            .I(II_1_counter_19));
    LocalMux I__555 (
            .O(N__2603),
            .I(II_1_counter_19));
    CascadeMux I__554 (
            .O(N__2594),
            .I(\II_1.un1_counterlto25_cascade_ ));
    InMux I__553 (
            .O(N__2591),
            .I(N__2584));
    InMux I__552 (
            .O(N__2590),
            .I(N__2581));
    InMux I__551 (
            .O(N__2589),
            .I(N__2576));
    InMux I__550 (
            .O(N__2588),
            .I(N__2576));
    InMux I__549 (
            .O(N__2587),
            .I(N__2573));
    LocalMux I__548 (
            .O(N__2584),
            .I(II_1_counter_18));
    LocalMux I__547 (
            .O(N__2581),
            .I(II_1_counter_18));
    LocalMux I__546 (
            .O(N__2576),
            .I(II_1_counter_18));
    LocalMux I__545 (
            .O(N__2573),
            .I(II_1_counter_18));
    InMux I__544 (
            .O(N__2564),
            .I(N__2561));
    LocalMux I__543 (
            .O(N__2561),
            .I(\II_1.counter_RNINVA12Z0Z_20 ));
    IoInMux I__542 (
            .O(N__2558),
            .I(N__2555));
    LocalMux I__541 (
            .O(N__2555),
            .I(N__2552));
    IoSpan4Mux I__540 (
            .O(N__2552),
            .I(N__2549));
    Span4Mux_s1_v I__539 (
            .O(N__2549),
            .I(N__2545));
    IoInMux I__538 (
            .O(N__2548),
            .I(N__2542));
    Span4Mux_h I__537 (
            .O(N__2545),
            .I(N__2535));
    LocalMux I__536 (
            .O(N__2542),
            .I(N__2535));
    IoInMux I__535 (
            .O(N__2541),
            .I(N__2531));
    InMux I__534 (
            .O(N__2540),
            .I(N__2528));
    Span4Mux_s1_v I__533 (
            .O(N__2535),
            .I(N__2525));
    IoInMux I__532 (
            .O(N__2534),
            .I(N__2522));
    LocalMux I__531 (
            .O(N__2531),
            .I(N__2519));
    LocalMux I__530 (
            .O(N__2528),
            .I(N__2516));
    Span4Mux_h I__529 (
            .O(N__2525),
            .I(N__2513));
    LocalMux I__528 (
            .O(N__2522),
            .I(N__2510));
    Span4Mux_s1_v I__527 (
            .O(N__2519),
            .I(N__2505));
    Span4Mux_v I__526 (
            .O(N__2516),
            .I(N__2505));
    Span4Mux_h I__525 (
            .O(N__2513),
            .I(N__2500));
    Span4Mux_s1_v I__524 (
            .O(N__2510),
            .I(N__2500));
    Sp12to4 I__523 (
            .O(N__2505),
            .I(N__2494));
    Sp12to4 I__522 (
            .O(N__2500),
            .I(N__2494));
    IoInMux I__521 (
            .O(N__2499),
            .I(N__2491));
    Span12Mux_h I__520 (
            .O(N__2494),
            .I(N__2488));
    LocalMux I__519 (
            .O(N__2491),
            .I(N__2485));
    Odrv12 I__518 (
            .O(N__2488),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__517 (
            .O(N__2485),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__516 (
            .O(N__2480),
            .I(\II_3.outputs_RNO_10Z0Z_0_cascade_ ));
    InMux I__515 (
            .O(N__2477),
            .I(N__2474));
    LocalMux I__514 (
            .O(N__2474),
            .I(N__2471));
    Odrv4 I__513 (
            .O(N__2471),
            .I(\II_3.G_30_0_a3_2_3 ));
    InMux I__512 (
            .O(N__2468),
            .I(N__2463));
    InMux I__511 (
            .O(N__2467),
            .I(N__2460));
    InMux I__510 (
            .O(N__2466),
            .I(N__2457));
    LocalMux I__509 (
            .O(N__2463),
            .I(\II_1.counterZ0Z_10 ));
    LocalMux I__508 (
            .O(N__2460),
            .I(\II_1.counterZ0Z_10 ));
    LocalMux I__507 (
            .O(N__2457),
            .I(\II_1.counterZ0Z_10 ));
    InMux I__506 (
            .O(N__2450),
            .I(N__2443));
    InMux I__505 (
            .O(N__2449),
            .I(N__2440));
    InMux I__504 (
            .O(N__2448),
            .I(N__2435));
    InMux I__503 (
            .O(N__2447),
            .I(N__2435));
    InMux I__502 (
            .O(N__2446),
            .I(N__2432));
    LocalMux I__501 (
            .O(N__2443),
            .I(II_1_counter_9));
    LocalMux I__500 (
            .O(N__2440),
            .I(II_1_counter_9));
    LocalMux I__499 (
            .O(N__2435),
            .I(II_1_counter_9));
    LocalMux I__498 (
            .O(N__2432),
            .I(II_1_counter_9));
    InMux I__497 (
            .O(N__2423),
            .I(N__2417));
    CascadeMux I__496 (
            .O(N__2422),
            .I(N__2413));
    InMux I__495 (
            .O(N__2421),
            .I(N__2410));
    InMux I__494 (
            .O(N__2420),
            .I(N__2407));
    LocalMux I__493 (
            .O(N__2417),
            .I(N__2404));
    InMux I__492 (
            .O(N__2416),
            .I(N__2401));
    InMux I__491 (
            .O(N__2413),
            .I(N__2398));
    LocalMux I__490 (
            .O(N__2410),
            .I(II_1_counter_11));
    LocalMux I__489 (
            .O(N__2407),
            .I(II_1_counter_11));
    Odrv4 I__488 (
            .O(N__2404),
            .I(II_1_counter_11));
    LocalMux I__487 (
            .O(N__2401),
            .I(II_1_counter_11));
    LocalMux I__486 (
            .O(N__2398),
            .I(II_1_counter_11));
    InMux I__485 (
            .O(N__2387),
            .I(N__2382));
    InMux I__484 (
            .O(N__2386),
            .I(N__2379));
    InMux I__483 (
            .O(N__2385),
            .I(N__2376));
    LocalMux I__482 (
            .O(N__2382),
            .I(\II_1.counterZ0Z_7 ));
    LocalMux I__481 (
            .O(N__2379),
            .I(\II_1.counterZ0Z_7 ));
    LocalMux I__480 (
            .O(N__2376),
            .I(\II_1.counterZ0Z_7 ));
    InMux I__479 (
            .O(N__2369),
            .I(N__2362));
    InMux I__478 (
            .O(N__2368),
            .I(N__2357));
    InMux I__477 (
            .O(N__2367),
            .I(N__2357));
    InMux I__476 (
            .O(N__2366),
            .I(N__2352));
    InMux I__475 (
            .O(N__2365),
            .I(N__2352));
    LocalMux I__474 (
            .O(N__2362),
            .I(II_1_counter_16));
    LocalMux I__473 (
            .O(N__2357),
            .I(II_1_counter_16));
    LocalMux I__472 (
            .O(N__2352),
            .I(II_1_counter_16));
    InMux I__471 (
            .O(N__2345),
            .I(N__2338));
    InMux I__470 (
            .O(N__2344),
            .I(N__2335));
    InMux I__469 (
            .O(N__2343),
            .I(N__2332));
    InMux I__468 (
            .O(N__2342),
            .I(N__2327));
    InMux I__467 (
            .O(N__2341),
            .I(N__2327));
    LocalMux I__466 (
            .O(N__2338),
            .I(II_1_counter_15));
    LocalMux I__465 (
            .O(N__2335),
            .I(II_1_counter_15));
    LocalMux I__464 (
            .O(N__2332),
            .I(II_1_counter_15));
    LocalMux I__463 (
            .O(N__2327),
            .I(II_1_counter_15));
    CascadeMux I__462 (
            .O(N__2318),
            .I(N__2311));
    InMux I__461 (
            .O(N__2317),
            .I(N__2308));
    InMux I__460 (
            .O(N__2316),
            .I(N__2303));
    InMux I__459 (
            .O(N__2315),
            .I(N__2303));
    InMux I__458 (
            .O(N__2314),
            .I(N__2298));
    InMux I__457 (
            .O(N__2311),
            .I(N__2298));
    LocalMux I__456 (
            .O(N__2308),
            .I(II_1_counter_17));
    LocalMux I__455 (
            .O(N__2303),
            .I(II_1_counter_17));
    LocalMux I__454 (
            .O(N__2298),
            .I(II_1_counter_17));
    InMux I__453 (
            .O(N__2291),
            .I(N__2287));
    InMux I__452 (
            .O(N__2290),
            .I(N__2281));
    LocalMux I__451 (
            .O(N__2287),
            .I(N__2278));
    InMux I__450 (
            .O(N__2286),
            .I(N__2271));
    InMux I__449 (
            .O(N__2285),
            .I(N__2271));
    InMux I__448 (
            .O(N__2284),
            .I(N__2271));
    LocalMux I__447 (
            .O(N__2281),
            .I(II_1_counter_14));
    Odrv4 I__446 (
            .O(N__2278),
            .I(II_1_counter_14));
    LocalMux I__445 (
            .O(N__2271),
            .I(II_1_counter_14));
    InMux I__444 (
            .O(N__2264),
            .I(N__2261));
    LocalMux I__443 (
            .O(N__2261),
            .I(N__2257));
    InMux I__442 (
            .O(N__2260),
            .I(N__2254));
    Span4Mux_s2_v I__441 (
            .O(N__2257),
            .I(N__2251));
    LocalMux I__440 (
            .O(N__2254),
            .I(\II_1.counterZ0Z_4 ));
    Odrv4 I__439 (
            .O(N__2251),
            .I(\II_1.counterZ0Z_4 ));
    CascadeMux I__438 (
            .O(N__2246),
            .I(N__2242));
    InMux I__437 (
            .O(N__2245),
            .I(N__2238));
    InMux I__436 (
            .O(N__2242),
            .I(N__2235));
    InMux I__435 (
            .O(N__2241),
            .I(N__2232));
    LocalMux I__434 (
            .O(N__2238),
            .I(N__2229));
    LocalMux I__433 (
            .O(N__2235),
            .I(N__2226));
    LocalMux I__432 (
            .O(N__2232),
            .I(\II_1.counterZ0Z_1 ));
    Odrv4 I__431 (
            .O(N__2229),
            .I(\II_1.counterZ0Z_1 ));
    Odrv4 I__430 (
            .O(N__2226),
            .I(\II_1.counterZ0Z_1 ));
    CascadeMux I__429 (
            .O(N__2219),
            .I(N__2216));
    InMux I__428 (
            .O(N__2216),
            .I(N__2212));
    InMux I__427 (
            .O(N__2215),
            .I(N__2209));
    LocalMux I__426 (
            .O(N__2212),
            .I(N__2206));
    LocalMux I__425 (
            .O(N__2209),
            .I(\II_1.counterZ0Z_5 ));
    Odrv4 I__424 (
            .O(N__2206),
            .I(\II_1.counterZ0Z_5 ));
    InMux I__423 (
            .O(N__2201),
            .I(N__2195));
    InMux I__422 (
            .O(N__2200),
            .I(N__2192));
    InMux I__421 (
            .O(N__2199),
            .I(N__2187));
    InMux I__420 (
            .O(N__2198),
            .I(N__2187));
    LocalMux I__419 (
            .O(N__2195),
            .I(N__2184));
    LocalMux I__418 (
            .O(N__2192),
            .I(N__2181));
    LocalMux I__417 (
            .O(N__2187),
            .I(\II_1.counterZ0Z_0 ));
    Odrv4 I__416 (
            .O(N__2184),
            .I(\II_1.counterZ0Z_0 ));
    Odrv4 I__415 (
            .O(N__2181),
            .I(\II_1.counterZ0Z_0 ));
    InMux I__414 (
            .O(N__2174),
            .I(N__2169));
    InMux I__413 (
            .O(N__2173),
            .I(N__2166));
    InMux I__412 (
            .O(N__2172),
            .I(N__2163));
    LocalMux I__411 (
            .O(N__2169),
            .I(\II_1.counterZ0Z_21 ));
    LocalMux I__410 (
            .O(N__2166),
            .I(\II_1.counterZ0Z_21 ));
    LocalMux I__409 (
            .O(N__2163),
            .I(\II_1.counterZ0Z_21 ));
    InMux I__408 (
            .O(N__2156),
            .I(N__2149));
    InMux I__407 (
            .O(N__2155),
            .I(N__2144));
    InMux I__406 (
            .O(N__2154),
            .I(N__2144));
    InMux I__405 (
            .O(N__2153),
            .I(N__2139));
    InMux I__404 (
            .O(N__2152),
            .I(N__2139));
    LocalMux I__403 (
            .O(N__2149),
            .I(II_1_counter_22));
    LocalMux I__402 (
            .O(N__2144),
            .I(II_1_counter_22));
    LocalMux I__401 (
            .O(N__2139),
            .I(II_1_counter_22));
    InMux I__400 (
            .O(N__2132),
            .I(N__2129));
    LocalMux I__399 (
            .O(N__2129),
            .I(N__2126));
    Odrv12 I__398 (
            .O(N__2126),
            .I(\II_1.un2_clock_outlto23_0_0_c ));
    CascadeMux I__397 (
            .O(N__2123),
            .I(N__2119));
    InMux I__396 (
            .O(N__2122),
            .I(N__2113));
    InMux I__395 (
            .O(N__2119),
            .I(N__2110));
    InMux I__394 (
            .O(N__2118),
            .I(N__2105));
    InMux I__393 (
            .O(N__2117),
            .I(N__2105));
    InMux I__392 (
            .O(N__2116),
            .I(N__2102));
    LocalMux I__391 (
            .O(N__2113),
            .I(II_1_counter_13));
    LocalMux I__390 (
            .O(N__2110),
            .I(II_1_counter_13));
    LocalMux I__389 (
            .O(N__2105),
            .I(II_1_counter_13));
    LocalMux I__388 (
            .O(N__2102),
            .I(II_1_counter_13));
    InMux I__387 (
            .O(N__2093),
            .I(N__2090));
    LocalMux I__386 (
            .O(N__2090),
            .I(\II_1.counter_RNIQ7FB1Z0Z_14 ));
    InMux I__385 (
            .O(N__2087),
            .I(N__2080));
    InMux I__384 (
            .O(N__2086),
            .I(N__2077));
    InMux I__383 (
            .O(N__2085),
            .I(N__2074));
    InMux I__382 (
            .O(N__2084),
            .I(N__2069));
    InMux I__381 (
            .O(N__2083),
            .I(N__2069));
    LocalMux I__380 (
            .O(N__2080),
            .I(N__2066));
    LocalMux I__379 (
            .O(N__2077),
            .I(II_1_counter_8));
    LocalMux I__378 (
            .O(N__2074),
            .I(II_1_counter_8));
    LocalMux I__377 (
            .O(N__2069),
            .I(II_1_counter_8));
    Odrv4 I__376 (
            .O(N__2066),
            .I(II_1_counter_8));
    CascadeMux I__375 (
            .O(N__2057),
            .I(\II_1.counter_RNI6VAM1Z0Z_13_cascade_ ));
    InMux I__374 (
            .O(N__2054),
            .I(N__2051));
    LocalMux I__373 (
            .O(N__2051),
            .I(\II_1.counter_RNIJ54VZ0Z_7 ));
    InMux I__372 (
            .O(N__2048),
            .I(bfn_15_32_0_));
    InMux I__371 (
            .O(N__2045),
            .I(\II_1.counter_1_cry_25 ));
    InMux I__370 (
            .O(N__2042),
            .I(\II_1.counter_1_cry_26 ));
    SRMux I__369 (
            .O(N__2039),
            .I(N__2024));
    SRMux I__368 (
            .O(N__2038),
            .I(N__2024));
    SRMux I__367 (
            .O(N__2037),
            .I(N__2024));
    SRMux I__366 (
            .O(N__2036),
            .I(N__2024));
    SRMux I__365 (
            .O(N__2035),
            .I(N__2024));
    GlobalMux I__364 (
            .O(N__2024),
            .I(N__2021));
    gio2CtrlBuf I__363 (
            .O(N__2021),
            .I(\II_1.un1_counter_0_g ));
    InMux I__362 (
            .O(N__2018),
            .I(N__2013));
    InMux I__361 (
            .O(N__2017),
            .I(N__2010));
    InMux I__360 (
            .O(N__2016),
            .I(N__2007));
    LocalMux I__359 (
            .O(N__2013),
            .I(\II_1.counterZ0Z_6 ));
    LocalMux I__358 (
            .O(N__2010),
            .I(\II_1.counterZ0Z_6 ));
    LocalMux I__357 (
            .O(N__2007),
            .I(\II_1.counterZ0Z_6 ));
    InMux I__356 (
            .O(N__2000),
            .I(N__1996));
    InMux I__355 (
            .O(N__1999),
            .I(N__1993));
    LocalMux I__354 (
            .O(N__1996),
            .I(\II_1.counterZ0Z_2 ));
    LocalMux I__353 (
            .O(N__1993),
            .I(\II_1.counterZ0Z_2 ));
    InMux I__352 (
            .O(N__1988),
            .I(N__1984));
    InMux I__351 (
            .O(N__1987),
            .I(N__1981));
    LocalMux I__350 (
            .O(N__1984),
            .I(\II_1.counterZ0Z_3 ));
    LocalMux I__349 (
            .O(N__1981),
            .I(\II_1.counterZ0Z_3 ));
    CascadeMux I__348 (
            .O(N__1976),
            .I(\II_1.un2_clock_outlto19_1_cascade_ ));
    InMux I__347 (
            .O(N__1973),
            .I(N__1970));
    LocalMux I__346 (
            .O(N__1970),
            .I(\II_1.un2_clock_outlto19_1 ));
    InMux I__345 (
            .O(N__1967),
            .I(N__1964));
    LocalMux I__344 (
            .O(N__1964),
            .I(N__1961));
    Span4Mux_h I__343 (
            .O(N__1961),
            .I(N__1958));
    Odrv4 I__342 (
            .O(N__1958),
            .I(\II_1.clock_out_RNOZ0Z_3 ));
    CascadeMux I__341 (
            .O(N__1955),
            .I(\II_1.un2_clock_outlto23_0_0_d_1_cascade_ ));
    InMux I__340 (
            .O(N__1952),
            .I(N__1949));
    LocalMux I__339 (
            .O(N__1949),
            .I(N__1945));
    InMux I__338 (
            .O(N__1948),
            .I(N__1942));
    Span4Mux_h I__337 (
            .O(N__1945),
            .I(N__1938));
    LocalMux I__336 (
            .O(N__1942),
            .I(N__1935));
    InMux I__335 (
            .O(N__1941),
            .I(N__1932));
    Odrv4 I__334 (
            .O(N__1938),
            .I(counter_RNIG1JB1_20));
    Odrv4 I__333 (
            .O(N__1935),
            .I(counter_RNIG1JB1_20));
    LocalMux I__332 (
            .O(N__1932),
            .I(counter_RNIG1JB1_20));
    CascadeMux I__331 (
            .O(N__1925),
            .I(\II_1.un2_clock_outlto23_0_0_d_cascade_ ));
    IoInMux I__330 (
            .O(N__1922),
            .I(N__1919));
    LocalMux I__329 (
            .O(N__1919),
            .I(N__1915));
    ClkMux I__328 (
            .O(N__1918),
            .I(N__1912));
    IoSpan4Mux I__327 (
            .O(N__1915),
            .I(N__1907));
    LocalMux I__326 (
            .O(N__1912),
            .I(N__1907));
    IoSpan4Mux I__325 (
            .O(N__1907),
            .I(N__1904));
    IoSpan4Mux I__324 (
            .O(N__1904),
            .I(N__1900));
    ClkMux I__323 (
            .O(N__1903),
            .I(N__1897));
    IoSpan4Mux I__322 (
            .O(N__1900),
            .I(N__1891));
    LocalMux I__321 (
            .O(N__1897),
            .I(N__1891));
    InMux I__320 (
            .O(N__1896),
            .I(N__1888));
    IoSpan4Mux I__319 (
            .O(N__1891),
            .I(N__1885));
    LocalMux I__318 (
            .O(N__1888),
            .I(N__1882));
    Span4Mux_s1_v I__317 (
            .O(N__1885),
            .I(N__1879));
    Span4Mux_s2_v I__316 (
            .O(N__1882),
            .I(N__1876));
    Odrv4 I__315 (
            .O(N__1879),
            .I(led8_c));
    Odrv4 I__314 (
            .O(N__1876),
            .I(led8_c));
    InMux I__313 (
            .O(N__1871),
            .I(N__1868));
    LocalMux I__312 (
            .O(N__1868),
            .I(N__1857));
    ClkMux I__311 (
            .O(N__1867),
            .I(N__1838));
    ClkMux I__310 (
            .O(N__1866),
            .I(N__1838));
    ClkMux I__309 (
            .O(N__1865),
            .I(N__1838));
    ClkMux I__308 (
            .O(N__1864),
            .I(N__1838));
    ClkMux I__307 (
            .O(N__1863),
            .I(N__1838));
    ClkMux I__306 (
            .O(N__1862),
            .I(N__1838));
    ClkMux I__305 (
            .O(N__1861),
            .I(N__1838));
    ClkMux I__304 (
            .O(N__1860),
            .I(N__1838));
    Glb2LocalMux I__303 (
            .O(N__1857),
            .I(N__1838));
    GlobalMux I__302 (
            .O(N__1838),
            .I(PLLOUTGLOBAL_0));
    InMux I__301 (
            .O(N__1835),
            .I(\II_1.counter_1_cry_15 ));
    InMux I__300 (
            .O(N__1832),
            .I(bfn_15_31_0_));
    InMux I__299 (
            .O(N__1829),
            .I(\II_1.counter_1_cry_17 ));
    InMux I__298 (
            .O(N__1826),
            .I(\II_1.counter_1_cry_18 ));
    InMux I__297 (
            .O(N__1823),
            .I(\II_1.counter_1_cry_19 ));
    InMux I__296 (
            .O(N__1820),
            .I(\II_1.counter_1_cry_20 ));
    InMux I__295 (
            .O(N__1817),
            .I(\II_1.counter_1_cry_21 ));
    InMux I__294 (
            .O(N__1814),
            .I(\II_1.counter_1_cry_22 ));
    InMux I__293 (
            .O(N__1811),
            .I(\II_1.counter_1_cry_23 ));
    InMux I__292 (
            .O(N__1808),
            .I(\II_1.counter_1_cry_6 ));
    InMux I__291 (
            .O(N__1805),
            .I(\II_1.counter_1_cry_7 ));
    InMux I__290 (
            .O(N__1802),
            .I(bfn_15_30_0_));
    InMux I__289 (
            .O(N__1799),
            .I(\II_1.counter_1_cry_9 ));
    InMux I__288 (
            .O(N__1796),
            .I(\II_1.counter_1_cry_10 ));
    InMux I__287 (
            .O(N__1793),
            .I(\II_1.counter_1_cry_11 ));
    InMux I__286 (
            .O(N__1790),
            .I(\II_1.counter_1_cry_12 ));
    InMux I__285 (
            .O(N__1787),
            .I(\II_1.counter_1_cry_13 ));
    InMux I__284 (
            .O(N__1784),
            .I(\II_1.counter_1_cry_14 ));
    InMux I__283 (
            .O(N__1781),
            .I(N__1778));
    LocalMux I__282 (
            .O(N__1778),
            .I(\II_3.G_30_0_o3_0 ));
    CascadeMux I__281 (
            .O(N__1775),
            .I(\II_1.counter_RNIM7JB1Z0Z_22_cascade_ ));
    InMux I__280 (
            .O(N__1772),
            .I(N__1769));
    LocalMux I__279 (
            .O(N__1769),
            .I(N__1766));
    Odrv4 I__278 (
            .O(N__1766),
            .I(\II_1.counter_RNI64GM1Z0Z_26 ));
    InMux I__277 (
            .O(N__1763),
            .I(\II_1.counter_1_cry_1 ));
    InMux I__276 (
            .O(N__1760),
            .I(\II_1.counter_1_cry_2 ));
    InMux I__275 (
            .O(N__1757),
            .I(\II_1.counter_1_cry_3 ));
    InMux I__274 (
            .O(N__1754),
            .I(\II_1.counter_1_cry_4 ));
    InMux I__273 (
            .O(N__1751),
            .I(\II_1.counter_1_cry_5 ));
    InMux I__272 (
            .O(N__1748),
            .I(N__1745));
    LocalMux I__271 (
            .O(N__1745),
            .I(\II_3.N_14 ));
    CascadeMux I__270 (
            .O(N__1742),
            .I(\II_3.G_30_0_o3_0_1_cascade_ ));
    InMux I__269 (
            .O(N__1739),
            .I(N__1736));
    LocalMux I__268 (
            .O(N__1736),
            .I(\II_1.counter_RNI1TC9Z0Z_8 ));
    InMux I__267 (
            .O(N__1733),
            .I(N__1730));
    LocalMux I__266 (
            .O(N__1730),
            .I(\II_3.N_16 ));
    InMux I__265 (
            .O(N__1727),
            .I(N__1724));
    LocalMux I__264 (
            .O(N__1724),
            .I(\II_3.G_30_0_a3_1 ));
    SRMux I__263 (
            .O(N__1721),
            .I(N__1718));
    LocalMux I__262 (
            .O(N__1718),
            .I(N__1715));
    Odrv4 I__261 (
            .O(N__1715),
            .I(\II_3.outputs_RNO_0Z0Z_0 ));
    CascadeMux I__260 (
            .O(N__1712),
            .I(N__1706));
    InMux I__259 (
            .O(N__1711),
            .I(N__1703));
    InMux I__258 (
            .O(N__1710),
            .I(N__1700));
    InMux I__257 (
            .O(N__1709),
            .I(N__1695));
    InMux I__256 (
            .O(N__1706),
            .I(N__1695));
    LocalMux I__255 (
            .O(N__1703),
            .I(N__1692));
    LocalMux I__254 (
            .O(N__1700),
            .I(N__1689));
    LocalMux I__253 (
            .O(N__1695),
            .I(\II_3.counterZ0Z_1 ));
    Odrv4 I__252 (
            .O(N__1692),
            .I(\II_3.counterZ0Z_1 ));
    Odrv4 I__251 (
            .O(N__1689),
            .I(\II_3.counterZ0Z_1 ));
    CascadeMux I__250 (
            .O(N__1682),
            .I(N__1678));
    InMux I__249 (
            .O(N__1681),
            .I(N__1674));
    InMux I__248 (
            .O(N__1678),
            .I(N__1670));
    InMux I__247 (
            .O(N__1677),
            .I(N__1667));
    LocalMux I__246 (
            .O(N__1674),
            .I(N__1664));
    InMux I__245 (
            .O(N__1673),
            .I(N__1661));
    LocalMux I__244 (
            .O(N__1670),
            .I(N__1656));
    LocalMux I__243 (
            .O(N__1667),
            .I(N__1656));
    Span4Mux_s1_v I__242 (
            .O(N__1664),
            .I(N__1653));
    LocalMux I__241 (
            .O(N__1661),
            .I(\II_3.counterZ0Z_2 ));
    Odrv4 I__240 (
            .O(N__1656),
            .I(\II_3.counterZ0Z_2 ));
    Odrv4 I__239 (
            .O(N__1653),
            .I(\II_3.counterZ0Z_2 ));
    InMux I__238 (
            .O(N__1646),
            .I(N__1639));
    InMux I__237 (
            .O(N__1645),
            .I(N__1636));
    InMux I__236 (
            .O(N__1644),
            .I(N__1629));
    InMux I__235 (
            .O(N__1643),
            .I(N__1629));
    InMux I__234 (
            .O(N__1642),
            .I(N__1629));
    LocalMux I__233 (
            .O(N__1639),
            .I(N__1626));
    LocalMux I__232 (
            .O(N__1636),
            .I(N__1623));
    LocalMux I__231 (
            .O(N__1629),
            .I(\II_3.counterZ0Z_0 ));
    Odrv4 I__230 (
            .O(N__1626),
            .I(\II_3.counterZ0Z_0 ));
    Odrv4 I__229 (
            .O(N__1623),
            .I(\II_3.counterZ0Z_0 ));
    CascadeMux I__228 (
            .O(N__1616),
            .I(\II_3.o2_0_cascade_ ));
    CascadeMux I__227 (
            .O(N__1613),
            .I(N__1610));
    InMux I__226 (
            .O(N__1610),
            .I(N__1607));
    LocalMux I__225 (
            .O(N__1607),
            .I(\II_3.N_12 ));
    InMux I__224 (
            .O(N__1604),
            .I(N__1580));
    InMux I__223 (
            .O(N__1603),
            .I(N__1580));
    InMux I__222 (
            .O(N__1602),
            .I(N__1580));
    InMux I__221 (
            .O(N__1601),
            .I(N__1580));
    InMux I__220 (
            .O(N__1600),
            .I(N__1580));
    InMux I__219 (
            .O(N__1599),
            .I(N__1580));
    InMux I__218 (
            .O(N__1598),
            .I(N__1580));
    InMux I__217 (
            .O(N__1597),
            .I(N__1580));
    LocalMux I__216 (
            .O(N__1580),
            .I(N__1574));
    InMux I__215 (
            .O(N__1579),
            .I(N__1571));
    InMux I__214 (
            .O(N__1578),
            .I(N__1568));
    InMux I__213 (
            .O(N__1577),
            .I(N__1565));
    Odrv4 I__212 (
            .O(N__1574),
            .I(II_2_G_3_out));
    LocalMux I__211 (
            .O(N__1571),
            .I(II_2_G_3_out));
    LocalMux I__210 (
            .O(N__1568),
            .I(II_2_G_3_out));
    LocalMux I__209 (
            .O(N__1565),
            .I(II_2_G_3_out));
    CascadeMux I__208 (
            .O(N__1556),
            .I(N__1550));
    CascadeMux I__207 (
            .O(N__1555),
            .I(N__1547));
    CascadeMux I__206 (
            .O(N__1554),
            .I(N__1544));
    InMux I__205 (
            .O(N__1553),
            .I(N__1533));
    InMux I__204 (
            .O(N__1550),
            .I(N__1533));
    InMux I__203 (
            .O(N__1547),
            .I(N__1533));
    InMux I__202 (
            .O(N__1544),
            .I(N__1533));
    InMux I__201 (
            .O(N__1543),
            .I(N__1530));
    InMux I__200 (
            .O(N__1542),
            .I(N__1527));
    LocalMux I__199 (
            .O(N__1533),
            .I(\II_2.counterZ0Z_2 ));
    LocalMux I__198 (
            .O(N__1530),
            .I(\II_2.counterZ0Z_2 ));
    LocalMux I__197 (
            .O(N__1527),
            .I(\II_2.counterZ0Z_2 ));
    CascadeMux I__196 (
            .O(N__1520),
            .I(N__1516));
    InMux I__195 (
            .O(N__1519),
            .I(N__1506));
    InMux I__194 (
            .O(N__1516),
            .I(N__1506));
    InMux I__193 (
            .O(N__1515),
            .I(N__1506));
    InMux I__192 (
            .O(N__1514),
            .I(N__1503));
    InMux I__191 (
            .O(N__1513),
            .I(N__1500));
    LocalMux I__190 (
            .O(N__1506),
            .I(\II_2.counterZ0Z_0 ));
    LocalMux I__189 (
            .O(N__1503),
            .I(\II_2.counterZ0Z_0 ));
    LocalMux I__188 (
            .O(N__1500),
            .I(\II_2.counterZ0Z_0 ));
    InMux I__187 (
            .O(N__1493),
            .I(N__1482));
    InMux I__186 (
            .O(N__1492),
            .I(N__1482));
    InMux I__185 (
            .O(N__1491),
            .I(N__1482));
    InMux I__184 (
            .O(N__1490),
            .I(N__1479));
    InMux I__183 (
            .O(N__1489),
            .I(N__1476));
    LocalMux I__182 (
            .O(N__1482),
            .I(\II_2.counterZ0Z_1 ));
    LocalMux I__181 (
            .O(N__1479),
            .I(\II_2.counterZ0Z_1 ));
    LocalMux I__180 (
            .O(N__1476),
            .I(\II_2.counterZ0Z_1 ));
    InMux I__179 (
            .O(N__1469),
            .I(N__1466));
    LocalMux I__178 (
            .O(N__1466),
            .I(\II_2.un1_counter19_1_0 ));
    CascadeMux I__177 (
            .O(N__1463),
            .I(counter_RNI6D8K_6_cascade_));
    InMux I__176 (
            .O(N__1460),
            .I(N__1456));
    InMux I__175 (
            .O(N__1459),
            .I(N__1453));
    LocalMux I__174 (
            .O(N__1456),
            .I(counter_RNI6D8K_6));
    LocalMux I__173 (
            .O(N__1453),
            .I(counter_RNI6D8K_6));
    CascadeMux I__172 (
            .O(N__1448),
            .I(\II_1.clock_out_RNOZ0Z_5_cascade_ ));
    InMux I__171 (
            .O(N__1445),
            .I(N__1442));
    LocalMux I__170 (
            .O(N__1442),
            .I(\II_1.counter_RNIK1FB1Z0Z_13 ));
    InMux I__169 (
            .O(N__1439),
            .I(N__1436));
    LocalMux I__168 (
            .O(N__1436),
            .I(\II_1.counter_RNIJLJ01_0Z0Z_17 ));
    InMux I__167 (
            .O(N__1433),
            .I(N__1430));
    LocalMux I__166 (
            .O(N__1430),
            .I(\II_1.un1_counterlt12_2 ));
    IoInMux I__165 (
            .O(N__1427),
            .I(N__1424));
    LocalMux I__164 (
            .O(N__1424),
            .I(N__1421));
    Span4Mux_s0_v I__163 (
            .O(N__1421),
            .I(N__1418));
    Span4Mux_h I__162 (
            .O(N__1418),
            .I(N__1415));
    Span4Mux_h I__161 (
            .O(N__1415),
            .I(N__1411));
    InMux I__160 (
            .O(N__1414),
            .I(N__1408));
    Odrv4 I__159 (
            .O(N__1411),
            .I(\II_2.outputsZ0Z_0 ));
    LocalMux I__158 (
            .O(N__1408),
            .I(\II_2.outputsZ0Z_0 ));
    CascadeMux I__157 (
            .O(N__1403),
            .I(\II_1.g3_3_cascade_ ));
    CascadeMux I__156 (
            .O(N__1400),
            .I(\II_1.counter_RNIIPRU2Z0Z_11_cascade_ ));
    InMux I__155 (
            .O(N__1397),
            .I(N__1394));
    LocalMux I__154 (
            .O(N__1394),
            .I(\II_1.g0_1_a4_0_0 ));
    CEMux I__153 (
            .O(N__1391),
            .I(N__1388));
    LocalMux I__152 (
            .O(N__1388),
            .I(N__1385));
    Span4Mux_v I__151 (
            .O(N__1385),
            .I(N__1381));
    InMux I__150 (
            .O(N__1384),
            .I(N__1378));
    Odrv4 I__149 (
            .O(N__1381),
            .I(II_1_un2_clock_outlt27_0_i));
    LocalMux I__148 (
            .O(N__1378),
            .I(II_1_un2_clock_outlt27_0_i));
    IoInMux I__147 (
            .O(N__1373),
            .I(N__1369));
    IoInMux I__146 (
            .O(N__1372),
            .I(N__1366));
    LocalMux I__145 (
            .O(N__1369),
            .I(N__1360));
    LocalMux I__144 (
            .O(N__1366),
            .I(N__1360));
    InMux I__143 (
            .O(N__1365),
            .I(N__1357));
    Odrv4 I__142 (
            .O(N__1360),
            .I(\II_3.outputsZ0Z_0 ));
    LocalMux I__141 (
            .O(N__1357),
            .I(\II_3.outputsZ0Z_0 ));
    CascadeMux I__140 (
            .O(N__1352),
            .I(\II_3.o2_cascade_ ));
    InMux I__139 (
            .O(N__1349),
            .I(N__1345));
    InMux I__138 (
            .O(N__1348),
            .I(N__1342));
    LocalMux I__137 (
            .O(N__1345),
            .I(\II_2.un1_counter23_1_5 ));
    LocalMux I__136 (
            .O(N__1342),
            .I(\II_2.un1_counter23_1_5 ));
    IoInMux I__135 (
            .O(N__1337),
            .I(N__1334));
    LocalMux I__134 (
            .O(N__1334),
            .I(N__1331));
    Span12Mux_s8_h I__133 (
            .O(N__1331),
            .I(N__1328));
    Odrv12 I__132 (
            .O(N__1328),
            .I(GB_BUFFER_PLLOUTGLOBAL_0_THRU_CO));
    IoInMux I__131 (
            .O(N__1325),
            .I(N__1322));
    LocalMux I__130 (
            .O(N__1322),
            .I(N__1319));
    IoSpan4Mux I__129 (
            .O(N__1319),
            .I(N__1316));
    Span4Mux_s0_v I__128 (
            .O(N__1316),
            .I(N__1312));
    CascadeMux I__127 (
            .O(N__1315),
            .I(N__1309));
    Span4Mux_h I__126 (
            .O(N__1312),
            .I(N__1306));
    InMux I__125 (
            .O(N__1309),
            .I(N__1303));
    Odrv4 I__124 (
            .O(N__1306),
            .I(\II_2.outputsZ0Z_1 ));
    LocalMux I__123 (
            .O(N__1303),
            .I(\II_2.outputsZ0Z_1 ));
    IoInMux I__122 (
            .O(N__1298),
            .I(N__1295));
    LocalMux I__121 (
            .O(N__1295),
            .I(N__1292));
    Span12Mux_s7_v I__120 (
            .O(N__1292),
            .I(N__1289));
    Span12Mux_h I__119 (
            .O(N__1289),
            .I(N__1286));
    Span12Mux_v I__118 (
            .O(N__1286),
            .I(N__1283));
    Odrv12 I__117 (
            .O(N__1283),
            .I(RESET_c));
    IoInMux I__116 (
            .O(N__1280),
            .I(N__1277));
    LocalMux I__115 (
            .O(N__1277),
            .I(N__1274));
    IoSpan4Mux I__114 (
            .O(N__1274),
            .I(N__1271));
    Span4Mux_s3_h I__113 (
            .O(N__1271),
            .I(N__1268));
    Sp12to4 I__112 (
            .O(N__1268),
            .I(N__1265));
    Span12Mux_v I__111 (
            .O(N__1265),
            .I(N__1262));
    Span12Mux_h I__110 (
            .O(N__1262),
            .I(N__1259));
    Odrv12 I__109 (
            .O(N__1259),
            .I(PLLOUTCORE_c));
    defparam IN_MUX_bfv_15_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_29_0_));
    defparam IN_MUX_bfv_15_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_30_0_ (
            .carryinitin(\II_1.counter_1_cry_8 ),
            .carryinitout(bfn_15_30_0_));
    defparam IN_MUX_bfv_15_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_31_0_ (
            .carryinitin(\II_1.counter_1_cry_16 ),
            .carryinitout(bfn_15_31_0_));
    defparam IN_MUX_bfv_15_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_32_0_ (
            .carryinitin(\II_1.counter_1_cry_24 ),
            .carryinitout(bfn_15_32_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \II_1.counter_RNIJGA99_0_27  (
            .USERSIGNALTOGLOBALBUFFER(N__2831),
            .GLOBALBUFFEROUTPUT(\II_1.un1_counter_0_g ));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam GB_BUFFER_PLLOUTGLOBAL_0_THRU_LUT4_0_LC_9_4_4.C_ON=1'b0;
    defparam GB_BUFFER_PLLOUTGLOBAL_0_THRU_LUT4_0_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PLLOUTGLOBAL_0_THRU_LUT4_0_LC_9_4_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_PLLOUTGLOBAL_0_THRU_LUT4_0_LC_9_4_4 (
            .in0(N__1871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_PLLOUTGLOBAL_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_2.counter_1_LC_13_29_0 .C_ON=1'b0;
    defparam \II_2.counter_1_LC_13_29_0 .SEQ_MODE=4'b1000;
    defparam \II_2.counter_1_LC_13_29_0 .LUT_INIT=16'b1101011110100000;
    LogicCell40 \II_2.counter_1_LC_13_29_0  (
            .in0(N__1598),
            .in1(N__1553),
            .in2(N__1520),
            .in3(N__1492),
            .lcout(\II_2.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_2.counter_0_LC_13_29_1 .C_ON=1'b0;
    defparam \II_2.counter_0_LC_13_29_1 .SEQ_MODE=4'b1000;
    defparam \II_2.counter_0_LC_13_29_1 .LUT_INIT=16'b1001001111001100;
    LogicCell40 \II_2.counter_0_LC_13_29_1  (
            .in0(N__1491),
            .in1(N__1515),
            .in2(N__1555),
            .in3(N__1597),
            .lcout(\II_2.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_2.outputs_1_LC_13_29_2 .C_ON=1'b0;
    defparam \II_2.outputs_1_LC_13_29_2 .SEQ_MODE=4'b1000;
    defparam \II_2.outputs_1_LC_13_29_2 .LUT_INIT=16'b1101000011110010;
    LogicCell40 \II_2.outputs_1_LC_13_29_2  (
            .in0(N__1601),
            .in1(N__1349),
            .in2(N__1315),
            .in3(N__1469),
            .lcout(\II_2.outputsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_2.counter_2_LC_13_29_3 .C_ON=1'b0;
    defparam \II_2.counter_2_LC_13_29_3 .SEQ_MODE=4'b1000;
    defparam \II_2.counter_2_LC_13_29_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \II_2.counter_2_LC_13_29_3  (
            .in0(N__1493),
            .in1(N__1519),
            .in2(N__1556),
            .in3(N__1599),
            .lcout(\II_2.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_3.counter_1_LC_13_29_4 .C_ON=1'b0;
    defparam \II_3.counter_1_LC_13_29_4 .SEQ_MODE=4'b1000;
    defparam \II_3.counter_1_LC_13_29_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \II_3.counter_1_LC_13_29_4  (
            .in0(N__1603),
            .in1(N__1643),
            .in2(_gnd_net_),
            .in3(N__1709),
            .lcout(\II_3.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_3.counter_2_LC_13_29_5 .C_ON=1'b0;
    defparam \II_3.counter_2_LC_13_29_5 .SEQ_MODE=4'b1000;
    defparam \II_3.counter_2_LC_13_29_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \II_3.counter_2_LC_13_29_5  (
            .in0(N__1644),
            .in1(N__1673),
            .in2(N__1712),
            .in3(N__1604),
            .lcout(\II_3.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_3.counter_0_LC_13_29_6 .C_ON=1'b0;
    defparam \II_3.counter_0_LC_13_29_6 .SEQ_MODE=4'b1000;
    defparam \II_3.counter_0_LC_13_29_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \II_3.counter_0_LC_13_29_6  (
            .in0(N__1602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1642),
            .lcout(\II_3.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_2.outputs_0_LC_13_29_7 .C_ON=1'b0;
    defparam \II_2.outputs_0_LC_13_29_7 .SEQ_MODE=4'b1000;
    defparam \II_2.outputs_0_LC_13_29_7 .LUT_INIT=16'b1000101110101010;
    LogicCell40 \II_2.outputs_0_LC_13_29_7  (
            .in0(N__1414),
            .in1(N__1348),
            .in2(N__1554),
            .in3(N__1600),
            .lcout(\II_2.outputsZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1863),
            .ce(N__1391),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIVSFM1_25_LC_13_30_1 .C_ON=1'b0;
    defparam \II_1.counter_RNIVSFM1_25_LC_13_30_1 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIVSFM1_25_LC_13_30_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \II_1.counter_RNIVSFM1_25_LC_13_30_1  (
            .in0(N__1941),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2779),
            .lcout(\II_1.g0_1_a4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNI1QAM1_14_LC_13_30_3 .C_ON=1'b0;
    defparam \II_1.counter_RNI1QAM1_14_LC_13_30_3 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNI1QAM1_14_LC_13_30_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \II_1.counter_RNI1QAM1_14_LC_13_30_3  (
            .in0(N__2540),
            .in1(N__1445),
            .in2(_gnd_net_),
            .in3(N__2291),
            .lcout(),
            .ltout(\II_1.g3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIIPRU2_11_LC_13_30_4 .C_ON=1'b0;
    defparam \II_1.counter_RNIIPRU2_11_LC_13_30_4 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIIPRU2_11_LC_13_30_4 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \II_1.counter_RNIIPRU2_11_LC_13_30_4  (
            .in0(N__1459),
            .in1(N__1739),
            .in2(N__1403),
            .in3(N__2423),
            .lcout(),
            .ltout(\II_1.counter_RNIIPRU2Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIAGFC7_11_LC_13_30_5 .C_ON=1'b0;
    defparam \II_1.counter_RNIAGFC7_11_LC_13_30_5 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIAGFC7_11_LC_13_30_5 .LUT_INIT=16'b1111101100110011;
    LogicCell40 \II_1.counter_RNIAGFC7_11_LC_13_30_5  (
            .in0(N__1439),
            .in1(N__1772),
            .in2(N__1400),
            .in3(N__1397),
            .lcout(II_1_un2_clock_outlt27_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_0_LC_13_31_0 .C_ON=1'b0;
    defparam \II_3.outputs_0_LC_13_31_0 .SEQ_MODE=4'b1001;
    defparam \II_3.outputs_0_LC_13_31_0 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \II_3.outputs_0_LC_13_31_0  (
            .in0(N__1365),
            .in1(N__1384),
            .in2(N__1682),
            .in3(N__1579),
            .lcout(\II_3.outputsZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1867),
            .ce(),
            .sr(N__1721));
    defparam \II_3.outputs_RNO_5_0_LC_13_32_0 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_5_0_LC_13_32_0 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_5_0_LC_13_32_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \II_3.outputs_RNO_5_0_LC_13_32_0  (
            .in0(N__2780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1710),
            .lcout(),
            .ltout(\II_3.o2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_1_0_LC_13_32_1 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_1_0_LC_13_32_1 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_1_0_LC_13_32_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \II_3.outputs_RNO_1_0_LC_13_32_1  (
            .in0(N__1677),
            .in1(N__1645),
            .in2(N__1352),
            .in3(N__1577),
            .lcout(\II_3.G_30_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_2.counter_RNIEL821_0_LC_14_28_5 .C_ON=1'b0;
    defparam \II_2.counter_RNIEL821_0_LC_14_28_5 .SEQ_MODE=4'b0000;
    defparam \II_2.counter_RNIEL821_0_LC_14_28_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \II_2.counter_RNIEL821_0_LC_14_28_5  (
            .in0(N__1542),
            .in1(N__1490),
            .in2(_gnd_net_),
            .in3(N__1514),
            .lcout(\II_2.un1_counter23_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_2.outputs_RNO_0_1_LC_14_29_0 .C_ON=1'b0;
    defparam \II_2.outputs_RNO_0_1_LC_14_29_0 .SEQ_MODE=4'b0000;
    defparam \II_2.outputs_RNO_0_1_LC_14_29_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \II_2.outputs_RNO_0_1_LC_14_29_0  (
            .in0(N__1543),
            .in1(N__1513),
            .in2(_gnd_net_),
            .in3(N__1489),
            .lcout(\II_2.un1_counter19_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNI6D8K_6_LC_14_29_1 .C_ON=1'b0;
    defparam \II_1.counter_RNI6D8K_6_LC_14_29_1 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNI6D8K_6_LC_14_29_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \II_1.counter_RNI6D8K_6_LC_14_29_1  (
            .in0(N__2017),
            .in1(N__2467),
            .in2(_gnd_net_),
            .in3(N__2386),
            .lcout(counter_RNI6D8K_6),
            .ltout(counter_RNI6D8K_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_9_0_LC_14_29_2 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_9_0_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_9_0_LC_14_29_2 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \II_3.outputs_RNO_9_0_LC_14_29_2  (
            .in0(N__2085),
            .in1(N__2416),
            .in2(N__1463),
            .in3(N__2449),
            .lcout(\II_3.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_RNO_5_LC_14_30_0 .C_ON=1'b0;
    defparam \II_1.clock_out_RNO_5_LC_14_30_0 .SEQ_MODE=4'b0000;
    defparam \II_1.clock_out_RNO_5_LC_14_30_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \II_1.clock_out_RNO_5_LC_14_30_0  (
            .in0(N__2118),
            .in1(N__2906),
            .in2(_gnd_net_),
            .in3(N__2368),
            .lcout(),
            .ltout(\II_1.clock_out_RNOZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_RNO_3_LC_14_30_1 .C_ON=1'b0;
    defparam \II_1.clock_out_RNO_3_LC_14_30_1 .SEQ_MODE=4'b0000;
    defparam \II_1.clock_out_RNO_3_LC_14_30_1 .LUT_INIT=16'b0111111100001111;
    LogicCell40 \II_1.clock_out_RNO_3_LC_14_30_1  (
            .in0(N__1433),
            .in1(N__1460),
            .in2(N__1448),
            .in3(N__2420),
            .lcout(\II_1.clock_out_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIK1FB1_13_LC_14_30_2 .C_ON=1'b0;
    defparam \II_1.counter_RNIK1FB1_13_LC_14_30_2 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIK1FB1_13_LC_14_30_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \II_1.counter_RNIK1FB1_13_LC_14_30_2  (
            .in0(N__2117),
            .in1(N__2367),
            .in2(N__2908),
            .in3(N__2343),
            .lcout(\II_1.counter_RNIK1FB1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIJLJ01_0_17_LC_14_30_3 .C_ON=1'b0;
    defparam \II_1.counter_RNIJLJ01_0_17_LC_14_30_3 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIJLJ01_0_17_LC_14_30_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \II_1.counter_RNIJLJ01_0_17_LC_14_30_3  (
            .in0(N__2619),
            .in1(N__2589),
            .in2(_gnd_net_),
            .in3(N__2316),
            .lcout(\II_1.counter_RNIJLJ01_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_RNO_4_LC_14_30_4 .C_ON=1'b0;
    defparam \II_1.clock_out_RNO_4_LC_14_30_4 .SEQ_MODE=4'b0000;
    defparam \II_1.clock_out_RNO_4_LC_14_30_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \II_1.clock_out_RNO_4_LC_14_30_4  (
            .in0(N__2084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2448),
            .lcout(\II_1.un1_counterlt12_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_8_0_LC_14_30_5 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_8_0_LC_14_30_5 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_8_0_LC_14_30_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \II_3.outputs_RNO_8_0_LC_14_30_5  (
            .in0(N__2618),
            .in1(N__2588),
            .in2(_gnd_net_),
            .in3(N__2315),
            .lcout(),
            .ltout(\II_3.G_30_0_o3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_4_0_LC_14_30_6 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_4_0_LC_14_30_6 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_4_0_LC_14_30_6 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \II_3.outputs_RNO_4_0_LC_14_30_6  (
            .in0(N__1748),
            .in1(N__1948),
            .in2(N__1742),
            .in3(N__2477),
            .lcout(\II_3.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNI1TC9_8_LC_14_30_7 .C_ON=1'b0;
    defparam \II_1.counter_RNI1TC9_8_LC_14_30_7 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNI1TC9_8_LC_14_30_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \II_1.counter_RNI1TC9_8_LC_14_30_7  (
            .in0(N__2447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2083),
            .lcout(\II_1.counter_RNI1TC9Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_1_LC_14_31_1 .C_ON=1'b0;
    defparam \II_1.counter_1_LC_14_31_1 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_1_LC_14_31_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \II_1.counter_1_LC_14_31_1  (
            .in0(N__2199),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2241),
            .lcout(\II_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1865),
            .ce(),
            .sr(N__2037));
    defparam \II_1.counter_RNIG1JB1_20_LC_14_31_2 .C_ON=1'b0;
    defparam \II_1.counter_RNIG1JB1_20_LC_14_31_2 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIG1JB1_20_LC_14_31_2 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \II_1.counter_RNIG1JB1_20_LC_14_31_2  (
            .in0(N__2716),
            .in1(N__2682),
            .in2(N__2645),
            .in3(N__2173),
            .lcout(counter_RNIG1JB1_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_0_LC_14_31_4 .C_ON=1'b0;
    defparam \II_1.counter_0_LC_14_31_4 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_0_LC_14_31_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \II_1.counter_0_LC_14_31_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2198),
            .lcout(\II_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1865),
            .ce(),
            .sr(N__2037));
    defparam \II_3.outputs_RNO_0_0_LC_14_31_6 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_0_0_LC_14_31_6 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_0_0_LC_14_31_6 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \II_3.outputs_RNO_0_0_LC_14_31_6  (
            .in0(N__1781),
            .in1(N__1733),
            .in2(N__1613),
            .in3(N__1727),
            .lcout(\II_3.outputs_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_6_0_LC_14_32_1 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_6_0_LC_14_32_1 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_6_0_LC_14_32_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \II_3.outputs_RNO_6_0_LC_14_32_1  (
            .in0(_gnd_net_),
            .in1(N__1711),
            .in2(_gnd_net_),
            .in3(N__2818),
            .lcout(),
            .ltout(\II_3.o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_3_0_LC_14_32_2 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_3_0_LC_14_32_2 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_3_0_LC_14_32_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \II_3.outputs_RNO_3_0_LC_14_32_2  (
            .in0(N__1681),
            .in1(N__1646),
            .in2(N__1616),
            .in3(N__1578),
            .lcout(\II_3.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_2.G_3_s_LC_14_32_3 .C_ON=1'b0;
    defparam \II_2.G_3_s_LC_14_32_3 .SEQ_MODE=4'b0000;
    defparam \II_2.G_3_s_LC_14_32_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \II_2.G_3_s_LC_14_32_3  (
            .in0(_gnd_net_),
            .in1(N__2855),
            .in2(_gnd_net_),
            .in3(N__1896),
            .lcout(II_2_G_3_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_2_0_LC_14_32_4 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_2_0_LC_14_32_4 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_2_0_LC_14_32_4 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \II_3.outputs_RNO_2_0_LC_14_32_4  (
            .in0(N__2718),
            .in1(N__2681),
            .in2(_gnd_net_),
            .in3(N__2155),
            .lcout(\II_3.G_30_0_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIM7JB1_22_LC_14_32_6 .C_ON=1'b0;
    defparam \II_1.counter_RNIM7JB1_22_LC_14_32_6 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIM7JB1_22_LC_14_32_6 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \II_1.counter_RNIM7JB1_22_LC_14_32_6  (
            .in0(N__2717),
            .in1(N__2680),
            .in2(N__2777),
            .in3(N__2154),
            .lcout(),
            .ltout(\II_1.counter_RNIM7JB1Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNI64GM1_26_LC_14_32_7 .C_ON=1'b0;
    defparam \II_1.counter_RNI64GM1_26_LC_14_32_7 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNI64GM1_26_LC_14_32_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \II_1.counter_RNI64GM1_26_LC_14_32_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1775),
            .in3(N__2819),
            .lcout(\II_1.counter_RNI64GM1Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_1_cry_1_c_LC_15_29_0 .C_ON=1'b1;
    defparam \II_1.counter_1_cry_1_c_LC_15_29_0 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_1_cry_1_c_LC_15_29_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \II_1.counter_1_cry_1_c_LC_15_29_0  (
            .in0(_gnd_net_),
            .in1(N__2201),
            .in2(N__2246),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_29_0_),
            .carryout(\II_1.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_2_LC_15_29_1 .C_ON=1'b1;
    defparam \II_1.counter_2_LC_15_29_1 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_2_LC_15_29_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_2_LC_15_29_1  (
            .in0(_gnd_net_),
            .in1(N__2000),
            .in2(_gnd_net_),
            .in3(N__1763),
            .lcout(\II_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_1 ),
            .carryout(\II_1.counter_1_cry_2 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_3_LC_15_29_2 .C_ON=1'b1;
    defparam \II_1.counter_3_LC_15_29_2 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_3_LC_15_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_3_LC_15_29_2  (
            .in0(_gnd_net_),
            .in1(N__1988),
            .in2(_gnd_net_),
            .in3(N__1760),
            .lcout(\II_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_2 ),
            .carryout(\II_1.counter_1_cry_3 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_4_LC_15_29_3 .C_ON=1'b1;
    defparam \II_1.counter_4_LC_15_29_3 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_4_LC_15_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_4_LC_15_29_3  (
            .in0(_gnd_net_),
            .in1(N__2260),
            .in2(_gnd_net_),
            .in3(N__1757),
            .lcout(\II_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_3 ),
            .carryout(\II_1.counter_1_cry_4 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_5_LC_15_29_4 .C_ON=1'b1;
    defparam \II_1.counter_5_LC_15_29_4 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_5_LC_15_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_5_LC_15_29_4  (
            .in0(_gnd_net_),
            .in1(N__2215),
            .in2(_gnd_net_),
            .in3(N__1754),
            .lcout(\II_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_4 ),
            .carryout(\II_1.counter_1_cry_5 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_6_LC_15_29_5 .C_ON=1'b1;
    defparam \II_1.counter_6_LC_15_29_5 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_6_LC_15_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_6_LC_15_29_5  (
            .in0(_gnd_net_),
            .in1(N__2018),
            .in2(_gnd_net_),
            .in3(N__1751),
            .lcout(\II_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_5 ),
            .carryout(\II_1.counter_1_cry_6 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_7_LC_15_29_6 .C_ON=1'b1;
    defparam \II_1.counter_7_LC_15_29_6 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_7_LC_15_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_7_LC_15_29_6  (
            .in0(_gnd_net_),
            .in1(N__2387),
            .in2(_gnd_net_),
            .in3(N__1808),
            .lcout(\II_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_6 ),
            .carryout(\II_1.counter_1_cry_7 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_8_LC_15_29_7 .C_ON=1'b1;
    defparam \II_1.counter_8_LC_15_29_7 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_8_LC_15_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_8_LC_15_29_7  (
            .in0(_gnd_net_),
            .in1(N__2086),
            .in2(_gnd_net_),
            .in3(N__1805),
            .lcout(II_1_counter_8),
            .ltout(),
            .carryin(\II_1.counter_1_cry_7 ),
            .carryout(\II_1.counter_1_cry_8 ),
            .clk(N__1861),
            .ce(),
            .sr(N__2039));
    defparam \II_1.counter_9_LC_15_30_0 .C_ON=1'b1;
    defparam \II_1.counter_9_LC_15_30_0 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_9_LC_15_30_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_9_LC_15_30_0  (
            .in0(_gnd_net_),
            .in1(N__2450),
            .in2(_gnd_net_),
            .in3(N__1802),
            .lcout(II_1_counter_9),
            .ltout(),
            .carryin(bfn_15_30_0_),
            .carryout(\II_1.counter_1_cry_9 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_10_LC_15_30_1 .C_ON=1'b1;
    defparam \II_1.counter_10_LC_15_30_1 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_10_LC_15_30_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_10_LC_15_30_1  (
            .in0(_gnd_net_),
            .in1(N__2468),
            .in2(_gnd_net_),
            .in3(N__1799),
            .lcout(\II_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_9 ),
            .carryout(\II_1.counter_1_cry_10 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_11_LC_15_30_2 .C_ON=1'b1;
    defparam \II_1.counter_11_LC_15_30_2 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_11_LC_15_30_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_11_LC_15_30_2  (
            .in0(_gnd_net_),
            .in1(N__2421),
            .in2(_gnd_net_),
            .in3(N__1796),
            .lcout(II_1_counter_11),
            .ltout(),
            .carryin(\II_1.counter_1_cry_10 ),
            .carryout(\II_1.counter_1_cry_11 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_12_LC_15_30_3 .C_ON=1'b1;
    defparam \II_1.counter_12_LC_15_30_3 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_12_LC_15_30_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_12_LC_15_30_3  (
            .in0(_gnd_net_),
            .in1(N__2907),
            .in2(_gnd_net_),
            .in3(N__1793),
            .lcout(II_1_counter_12),
            .ltout(),
            .carryin(\II_1.counter_1_cry_11 ),
            .carryout(\II_1.counter_1_cry_12 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_13_LC_15_30_4 .C_ON=1'b1;
    defparam \II_1.counter_13_LC_15_30_4 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_13_LC_15_30_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_13_LC_15_30_4  (
            .in0(_gnd_net_),
            .in1(N__2122),
            .in2(_gnd_net_),
            .in3(N__1790),
            .lcout(II_1_counter_13),
            .ltout(),
            .carryin(\II_1.counter_1_cry_12 ),
            .carryout(\II_1.counter_1_cry_13 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_14_LC_15_30_5 .C_ON=1'b1;
    defparam \II_1.counter_14_LC_15_30_5 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_14_LC_15_30_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_14_LC_15_30_5  (
            .in0(_gnd_net_),
            .in1(N__2290),
            .in2(_gnd_net_),
            .in3(N__1787),
            .lcout(II_1_counter_14),
            .ltout(),
            .carryin(\II_1.counter_1_cry_13 ),
            .carryout(\II_1.counter_1_cry_14 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_15_LC_15_30_6 .C_ON=1'b1;
    defparam \II_1.counter_15_LC_15_30_6 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_15_LC_15_30_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_15_LC_15_30_6  (
            .in0(_gnd_net_),
            .in1(N__2345),
            .in2(_gnd_net_),
            .in3(N__1784),
            .lcout(II_1_counter_15),
            .ltout(),
            .carryin(\II_1.counter_1_cry_14 ),
            .carryout(\II_1.counter_1_cry_15 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_16_LC_15_30_7 .C_ON=1'b1;
    defparam \II_1.counter_16_LC_15_30_7 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_16_LC_15_30_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_16_LC_15_30_7  (
            .in0(_gnd_net_),
            .in1(N__2369),
            .in2(_gnd_net_),
            .in3(N__1835),
            .lcout(II_1_counter_16),
            .ltout(),
            .carryin(\II_1.counter_1_cry_15 ),
            .carryout(\II_1.counter_1_cry_16 ),
            .clk(N__1862),
            .ce(),
            .sr(N__2038));
    defparam \II_1.counter_17_LC_15_31_0 .C_ON=1'b1;
    defparam \II_1.counter_17_LC_15_31_0 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_17_LC_15_31_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_17_LC_15_31_0  (
            .in0(_gnd_net_),
            .in1(N__2317),
            .in2(_gnd_net_),
            .in3(N__1832),
            .lcout(II_1_counter_17),
            .ltout(),
            .carryin(bfn_15_31_0_),
            .carryout(\II_1.counter_1_cry_17 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_18_LC_15_31_1 .C_ON=1'b1;
    defparam \II_1.counter_18_LC_15_31_1 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_18_LC_15_31_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_18_LC_15_31_1  (
            .in0(_gnd_net_),
            .in1(N__2591),
            .in2(_gnd_net_),
            .in3(N__1829),
            .lcout(II_1_counter_18),
            .ltout(),
            .carryin(\II_1.counter_1_cry_17 ),
            .carryout(\II_1.counter_1_cry_18 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_19_LC_15_31_2 .C_ON=1'b1;
    defparam \II_1.counter_19_LC_15_31_2 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_19_LC_15_31_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_19_LC_15_31_2  (
            .in0(_gnd_net_),
            .in1(N__2621),
            .in2(_gnd_net_),
            .in3(N__1826),
            .lcout(II_1_counter_19),
            .ltout(),
            .carryin(\II_1.counter_1_cry_18 ),
            .carryout(\II_1.counter_1_cry_19 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_20_LC_15_31_3 .C_ON=1'b1;
    defparam \II_1.counter_20_LC_15_31_3 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_20_LC_15_31_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_20_LC_15_31_3  (
            .in0(_gnd_net_),
            .in1(N__2643),
            .in2(_gnd_net_),
            .in3(N__1823),
            .lcout(\II_1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_19 ),
            .carryout(\II_1.counter_1_cry_20 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_21_LC_15_31_4 .C_ON=1'b1;
    defparam \II_1.counter_21_LC_15_31_4 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_21_LC_15_31_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_21_LC_15_31_4  (
            .in0(_gnd_net_),
            .in1(N__2174),
            .in2(_gnd_net_),
            .in3(N__1820),
            .lcout(\II_1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\II_1.counter_1_cry_20 ),
            .carryout(\II_1.counter_1_cry_21 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_22_LC_15_31_5 .C_ON=1'b1;
    defparam \II_1.counter_22_LC_15_31_5 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_22_LC_15_31_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_22_LC_15_31_5  (
            .in0(_gnd_net_),
            .in1(N__2156),
            .in2(_gnd_net_),
            .in3(N__1817),
            .lcout(II_1_counter_22),
            .ltout(),
            .carryin(\II_1.counter_1_cry_21 ),
            .carryout(\II_1.counter_1_cry_22 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_23_LC_15_31_6 .C_ON=1'b1;
    defparam \II_1.counter_23_LC_15_31_6 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_23_LC_15_31_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_23_LC_15_31_6  (
            .in0(_gnd_net_),
            .in1(N__2683),
            .in2(_gnd_net_),
            .in3(N__1814),
            .lcout(II_1_counter_23),
            .ltout(),
            .carryin(\II_1.counter_1_cry_22 ),
            .carryout(\II_1.counter_1_cry_23 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_24_LC_15_31_7 .C_ON=1'b1;
    defparam \II_1.counter_24_LC_15_31_7 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_24_LC_15_31_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_24_LC_15_31_7  (
            .in0(_gnd_net_),
            .in1(N__2722),
            .in2(_gnd_net_),
            .in3(N__1811),
            .lcout(II_1_counter_24),
            .ltout(),
            .carryin(\II_1.counter_1_cry_23 ),
            .carryout(\II_1.counter_1_cry_24 ),
            .clk(N__1864),
            .ce(),
            .sr(N__2036));
    defparam \II_1.counter_25_LC_15_32_0 .C_ON=1'b1;
    defparam \II_1.counter_25_LC_15_32_0 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_25_LC_15_32_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_25_LC_15_32_0  (
            .in0(_gnd_net_),
            .in1(N__2769),
            .in2(_gnd_net_),
            .in3(N__2048),
            .lcout(II_1_counter_25),
            .ltout(),
            .carryin(bfn_15_32_0_),
            .carryout(\II_1.counter_1_cry_25 ),
            .clk(N__1866),
            .ce(),
            .sr(N__2035));
    defparam \II_1.counter_26_LC_15_32_1 .C_ON=1'b1;
    defparam \II_1.counter_26_LC_15_32_1 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_26_LC_15_32_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \II_1.counter_26_LC_15_32_1  (
            .in0(_gnd_net_),
            .in1(N__2820),
            .in2(_gnd_net_),
            .in3(N__2045),
            .lcout(II_1_counter_26),
            .ltout(),
            .carryin(\II_1.counter_1_cry_25 ),
            .carryout(\II_1.counter_1_cry_26 ),
            .clk(N__1866),
            .ce(),
            .sr(N__2035));
    defparam \II_1.counter_27_LC_15_32_2 .C_ON=1'b0;
    defparam \II_1.counter_27_LC_15_32_2 .SEQ_MODE=4'b1000;
    defparam \II_1.counter_27_LC_15_32_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \II_1.counter_27_LC_15_32_2  (
            .in0(_gnd_net_),
            .in1(N__2860),
            .in2(_gnd_net_),
            .in3(N__2042),
            .lcout(II_1_counter_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1866),
            .ce(),
            .sr(N__2035));
    defparam \II_1.counter_RNIJS2E_2_LC_16_29_0 .C_ON=1'b0;
    defparam \II_1.counter_RNIJS2E_2_LC_16_29_0 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIJS2E_2_LC_16_29_0 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \II_1.counter_RNIJS2E_2_LC_16_29_0  (
            .in0(N__2016),
            .in1(N__1999),
            .in2(_gnd_net_),
            .in3(N__1987),
            .lcout(\II_1.counter_RNIJS2EZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIJLJ01_17_LC_16_30_0 .C_ON=1'b0;
    defparam \II_1.counter_RNIJLJ01_17_LC_16_30_0 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIJLJ01_17_LC_16_30_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \II_1.counter_RNIJLJ01_17_LC_16_30_0  (
            .in0(N__2590),
            .in1(N__2620),
            .in2(_gnd_net_),
            .in3(N__2314),
            .lcout(\II_1.un2_clock_outlto19_1 ),
            .ltout(\II_1.un2_clock_outlto19_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_RNO_2_LC_16_30_1 .C_ON=1'b0;
    defparam \II_1.clock_out_RNO_2_LC_16_30_1 .SEQ_MODE=4'b0000;
    defparam \II_1.clock_out_RNO_2_LC_16_30_1 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \II_1.clock_out_RNO_2_LC_16_30_1  (
            .in0(N__2778),
            .in1(N__2342),
            .in2(N__1976),
            .in3(N__2286),
            .lcout(),
            .ltout(\II_1.un2_clock_outlto23_0_0_d_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_RNO_1_LC_16_30_2 .C_ON=1'b0;
    defparam \II_1.clock_out_RNO_1_LC_16_30_2 .SEQ_MODE=4'b0000;
    defparam \II_1.clock_out_RNO_1_LC_16_30_2 .LUT_INIT=16'b1000111111111111;
    LogicCell40 \II_1.clock_out_RNO_1_LC_16_30_2  (
            .in0(N__1973),
            .in1(N__1967),
            .in2(N__1955),
            .in3(N__1952),
            .lcout(),
            .ltout(\II_1.un2_clock_outlto23_0_0_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_LC_16_30_3 .C_ON=1'b0;
    defparam \II_1.clock_out_LC_16_30_3 .SEQ_MODE=4'b1000;
    defparam \II_1.clock_out_LC_16_30_3 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \II_1.clock_out_LC_16_30_3  (
            .in0(N__2132),
            .in1(N__2861),
            .in2(N__1925),
            .in3(N__2825),
            .lcout(led8_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1860),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_10_0_LC_16_30_4 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_10_0_LC_16_30_4 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_10_0_LC_16_30_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \II_3.outputs_RNO_10_0_LC_16_30_4  (
            .in0(N__2285),
            .in1(N__2366),
            .in2(N__2123),
            .in3(N__2344),
            .lcout(),
            .ltout(\II_3.outputs_RNO_10Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_3.outputs_RNO_7_0_LC_16_30_5 .C_ON=1'b0;
    defparam \II_3.outputs_RNO_7_0_LC_16_30_5 .SEQ_MODE=4'b0000;
    defparam \II_3.outputs_RNO_7_0_LC_16_30_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \II_3.outputs_RNO_7_0_LC_16_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2480),
            .in3(N__2905),
            .lcout(\II_3.G_30_0_a3_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIJ54V_7_LC_16_30_6 .C_ON=1'b0;
    defparam \II_1.counter_RNIJ54V_7_LC_16_30_6 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIJ54V_7_LC_16_30_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \II_1.counter_RNIJ54V_7_LC_16_30_6  (
            .in0(N__2466),
            .in1(N__2446),
            .in2(N__2422),
            .in3(N__2385),
            .lcout(\II_1.counter_RNIJ54VZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIQ7FB1_14_LC_16_30_7 .C_ON=1'b0;
    defparam \II_1.counter_RNIQ7FB1_14_LC_16_30_7 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIQ7FB1_14_LC_16_30_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \II_1.counter_RNIQ7FB1_14_LC_16_30_7  (
            .in0(N__2365),
            .in1(N__2341),
            .in2(N__2318),
            .in3(N__2284),
            .lcout(\II_1.counter_RNIQ7FB1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIA1PI_1_LC_16_31_0 .C_ON=1'b0;
    defparam \II_1.counter_RNIA1PI_1_LC_16_31_0 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIA1PI_1_LC_16_31_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \II_1.counter_RNIA1PI_1_LC_16_31_0  (
            .in0(N__2264),
            .in1(N__2245),
            .in2(N__2219),
            .in3(N__2200),
            .lcout(\II_1.counter_RNIA1PIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNINFPL_21_LC_16_31_3 .C_ON=1'b0;
    defparam \II_1.counter_RNINFPL_21_LC_16_31_3 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNINFPL_21_LC_16_31_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \II_1.counter_RNINFPL_21_LC_16_31_3  (
            .in0(_gnd_net_),
            .in1(N__2152),
            .in2(_gnd_net_),
            .in3(N__2172),
            .lcout(\II_1.un1_counterlto22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.clock_out_RNO_0_LC_16_31_5 .C_ON=1'b0;
    defparam \II_1.clock_out_RNO_0_LC_16_31_5 .SEQ_MODE=4'b0000;
    defparam \II_1.clock_out_RNO_0_LC_16_31_5 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \II_1.clock_out_RNO_0_LC_16_31_5  (
            .in0(N__2684),
            .in1(N__2765),
            .in2(N__2726),
            .in3(N__2153),
            .lcout(\II_1.un2_clock_outlto23_0_0_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNI6VAM1_13_LC_16_31_6 .C_ON=1'b0;
    defparam \II_1.counter_RNI6VAM1_13_LC_16_31_6 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNI6VAM1_13_LC_16_31_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \II_1.counter_RNI6VAM1_13_LC_16_31_6  (
            .in0(_gnd_net_),
            .in1(N__2116),
            .in2(_gnd_net_),
            .in3(N__2093),
            .lcout(),
            .ltout(\II_1.counter_RNI6VAM1Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNI49153_8_LC_16_31_7 .C_ON=1'b0;
    defparam \II_1.counter_RNI49153_8_LC_16_31_7 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNI49153_8_LC_16_31_7 .LUT_INIT=16'b0000010100100101;
    LogicCell40 \II_1.counter_RNI49153_8_LC_16_31_7  (
            .in0(N__2901),
            .in1(N__2087),
            .in2(N__2057),
            .in3(N__2054),
            .lcout(\II_1.counter_RNI49153Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNICTOG4_12_LC_16_32_0 .C_ON=1'b0;
    defparam \II_1.counter_RNICTOG4_12_LC_16_32_0 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNICTOG4_12_LC_16_32_0 .LUT_INIT=16'b1110000000001111;
    LogicCell40 \II_1.counter_RNICTOG4_12_LC_16_32_0  (
            .in0(N__2927),
            .in1(N__2921),
            .in2(N__2912),
            .in3(N__2867),
            .lcout(),
            .ltout(\II_1.counter_RNICTOG4Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIJGA99_27_LC_16_32_1 .C_ON=1'b0;
    defparam \II_1.counter_RNIJGA99_27_LC_16_32_1 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIJGA99_27_LC_16_32_1 .LUT_INIT=16'b0000100010101010;
    LogicCell40 \II_1.counter_RNIJGA99_27_LC_16_32_1  (
            .in0(N__2856),
            .in1(N__2564),
            .in2(N__2834),
            .in3(N__2786),
            .lcout(\II_1.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIVL9C2_26_LC_16_32_5 .C_ON=1'b0;
    defparam \II_1.counter_RNIVL9C2_26_LC_16_32_5 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIVL9C2_26_LC_16_32_5 .LUT_INIT=16'b0000011100000011;
    LogicCell40 \II_1.counter_RNIVL9C2_26_LC_16_32_5  (
            .in0(N__2715),
            .in1(N__2651),
            .in2(N__2824),
            .in3(N__2792),
            .lcout(\II_1.un1_counterlto24_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNIAFM01_23_LC_16_32_6 .C_ON=1'b0;
    defparam \II_1.counter_RNIAFM01_23_LC_16_32_6 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNIAFM01_23_LC_16_32_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \II_1.counter_RNIAFM01_23_LC_16_32_6  (
            .in0(N__2770),
            .in1(N__2714),
            .in2(_gnd_net_),
            .in3(N__2679),
            .lcout(\II_1.un1_counterlto25 ),
            .ltout(\II_1.un1_counterlto25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \II_1.counter_RNINVA12_20_LC_16_32_7 .C_ON=1'b0;
    defparam \II_1.counter_RNINVA12_20_LC_16_32_7 .SEQ_MODE=4'b0000;
    defparam \II_1.counter_RNINVA12_20_LC_16_32_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \II_1.counter_RNINVA12_20_LC_16_32_7  (
            .in0(N__2644),
            .in1(N__2617),
            .in2(N__2594),
            .in3(N__2587),
            .lcout(\II_1.counter_RNINVA12Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_27_31_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_27_31_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_27_31_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_27_31_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top_pll
