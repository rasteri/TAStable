-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Nov 8 2023 16:58:30

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top_pll" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top_pll
entity top_pll is
port (
    led6 : out std_logic;
    led2 : out std_logic;
    lcol1 : out std_logic;
    RESET : in std_logic;
    led7 : out std_logic;
    led3 : out std_logic;
    lcol4 : out std_logic;
    PLLOUTCORE : out std_logic;
    PACKAGEPIN : in std_logic;
    led8 : out std_logic;
    led4 : out std_logic;
    lcol3 : out std_logic;
    led5 : out std_logic;
    led1 : out std_logic;
    lcol2 : out std_logic;
    PLLOUTGLOBAL : out std_logic);
end top_pll;

-- Architecture of top_pll
-- View name is \INTERFACE\
architecture \INTERFACE\ of top_pll is

signal \N__3086\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2013\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1888\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1865\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1790\ : std_logic;
signal \N__1787\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1772\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1754\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1748\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1733\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1727\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1711\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1674\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1644\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1636\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1565\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1554\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1491\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1479\ : std_logic;
signal \N__1476\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1459\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1414\ : std_logic;
signal \N__1411\ : std_logic;
signal \N__1408\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1384\ : std_logic;
signal \N__1381\ : std_logic;
signal \N__1378\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1372\ : std_logic;
signal \N__1369\ : std_logic;
signal \N__1366\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1360\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1352\ : std_logic;
signal \N__1349\ : std_logic;
signal \N__1348\ : std_logic;
signal \N__1345\ : std_logic;
signal \N__1342\ : std_logic;
signal \N__1337\ : std_logic;
signal \N__1334\ : std_logic;
signal \N__1331\ : std_logic;
signal \N__1328\ : std_logic;
signal \N__1325\ : std_logic;
signal \N__1322\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1312\ : std_logic;
signal \N__1309\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1303\ : std_logic;
signal \N__1298\ : std_logic;
signal \N__1295\ : std_logic;
signal \N__1292\ : std_logic;
signal \N__1289\ : std_logic;
signal \N__1286\ : std_logic;
signal \N__1283\ : std_logic;
signal \N__1280\ : std_logic;
signal \N__1277\ : std_logic;
signal \N__1274\ : std_logic;
signal \N__1271\ : std_logic;
signal \N__1268\ : std_logic;
signal \N__1265\ : std_logic;
signal \N__1262\ : std_logic;
signal \N__1259\ : std_logic;
signal \VCCG0\ : std_logic;
signal \RESET_c\ : std_logic;
signal \PLLOUTCORE_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \GB_BUFFER_PLLOUTGLOBAL_0_THRU_CO\ : std_logic;
signal \II_2.outputsZ0Z_1\ : std_logic;
signal \II_2.outputsZ0Z_0\ : std_logic;
signal \II_1.g3_3_cascade_\ : std_logic;
signal \II_1.counter_RNIIPRU2Z0Z_11_cascade_\ : std_logic;
signal \II_1.g0_1_a4_0_0\ : std_logic;
signal \II_1_un2_clock_outlt27_0_i\ : std_logic;
signal \II_3.outputsZ0Z_0\ : std_logic;
signal \II_3.o2_cascade_\ : std_logic;
signal \II_2.un1_counter23_1_5\ : std_logic;
signal \II_2.counterZ0Z_2\ : std_logic;
signal \II_2.counterZ0Z_0\ : std_logic;
signal \II_2.counterZ0Z_1\ : std_logic;
signal \II_2.un1_counter19_1_0\ : std_logic;
signal \counter_RNI6D8K_6_cascade_\ : std_logic;
signal \counter_RNI6D8K_6\ : std_logic;
signal \II_1.clock_out_RNOZ0Z_5_cascade_\ : std_logic;
signal \II_1.counter_RNIK1FB1Z0Z_13\ : std_logic;
signal \II_1.counter_RNIJLJ01_0Z0Z_17\ : std_logic;
signal \II_1.un1_counterlt12_2\ : std_logic;
signal \II_3.N_14\ : std_logic;
signal \II_3.G_30_0_o3_0_1_cascade_\ : std_logic;
signal \II_1.counter_RNI1TC9Z0Z_8\ : std_logic;
signal \II_3.N_16\ : std_logic;
signal \II_3.G_30_0_a3_1\ : std_logic;
signal \II_3.outputs_RNO_0Z0Z_0\ : std_logic;
signal \II_3.counterZ0Z_1\ : std_logic;
signal \II_3.counterZ0Z_2\ : std_logic;
signal \II_3.counterZ0Z_0\ : std_logic;
signal \II_3.o2_0_cascade_\ : std_logic;
signal \II_3.N_12\ : std_logic;
signal \II_2_G_3_out\ : std_logic;
signal \II_3.G_30_0_o3_0\ : std_logic;
signal \II_1.counter_RNIM7JB1Z0Z_22_cascade_\ : std_logic;
signal \II_1.counter_RNI64GM1Z0Z_26\ : std_logic;
signal \bfn_15_29_0_\ : std_logic;
signal \II_1.counter_1_cry_1\ : std_logic;
signal \II_1.counter_1_cry_2\ : std_logic;
signal \II_1.counter_1_cry_3\ : std_logic;
signal \II_1.counter_1_cry_4\ : std_logic;
signal \II_1.counter_1_cry_5\ : std_logic;
signal \II_1.counter_1_cry_6\ : std_logic;
signal \II_1.counter_1_cry_7\ : std_logic;
signal \II_1.counter_1_cry_8\ : std_logic;
signal \bfn_15_30_0_\ : std_logic;
signal \II_1.counter_1_cry_9\ : std_logic;
signal \II_1.counter_1_cry_10\ : std_logic;
signal \II_1.counter_1_cry_11\ : std_logic;
signal \II_1.counter_1_cry_12\ : std_logic;
signal \II_1.counter_1_cry_13\ : std_logic;
signal \II_1.counter_1_cry_14\ : std_logic;
signal \II_1.counter_1_cry_15\ : std_logic;
signal \II_1.counter_1_cry_16\ : std_logic;
signal \bfn_15_31_0_\ : std_logic;
signal \II_1.counter_1_cry_17\ : std_logic;
signal \II_1.counter_1_cry_18\ : std_logic;
signal \II_1.counter_1_cry_19\ : std_logic;
signal \II_1.counter_1_cry_20\ : std_logic;
signal \II_1.counter_1_cry_21\ : std_logic;
signal \II_1.counter_1_cry_22\ : std_logic;
signal \II_1.counter_1_cry_23\ : std_logic;
signal \II_1.counter_1_cry_24\ : std_logic;
signal \bfn_15_32_0_\ : std_logic;
signal \II_1.counter_1_cry_25\ : std_logic;
signal \II_1.counter_1_cry_26\ : std_logic;
signal \II_1.un1_counter_0_g\ : std_logic;
signal \II_1.counterZ0Z_6\ : std_logic;
signal \II_1.counterZ0Z_2\ : std_logic;
signal \II_1.counterZ0Z_3\ : std_logic;
signal \II_1.un2_clock_outlto19_1_cascade_\ : std_logic;
signal \II_1.un2_clock_outlto19_1\ : std_logic;
signal \II_1.clock_out_RNOZ0Z_3\ : std_logic;
signal \II_1.un2_clock_outlto23_0_0_d_1_cascade_\ : std_logic;
signal \counter_RNIG1JB1_20\ : std_logic;
signal \II_1.un2_clock_outlto23_0_0_d_cascade_\ : std_logic;
signal led8_c : std_logic;
signal \PLLOUTGLOBAL_0\ : std_logic;
signal \II_3.outputs_RNO_10Z0Z_0_cascade_\ : std_logic;
signal \II_3.G_30_0_a3_2_3\ : std_logic;
signal \II_1.counterZ0Z_10\ : std_logic;
signal \II_1_counter_9\ : std_logic;
signal \II_1_counter_11\ : std_logic;
signal \II_1.counterZ0Z_7\ : std_logic;
signal \II_1_counter_16\ : std_logic;
signal \II_1_counter_15\ : std_logic;
signal \II_1_counter_17\ : std_logic;
signal \II_1_counter_14\ : std_logic;
signal \II_1.counterZ0Z_4\ : std_logic;
signal \II_1.counterZ0Z_1\ : std_logic;
signal \II_1.counterZ0Z_5\ : std_logic;
signal \II_1.counterZ0Z_0\ : std_logic;
signal \II_1.counterZ0Z_21\ : std_logic;
signal \II_1_counter_22\ : std_logic;
signal \II_1.un2_clock_outlto23_0_0_c\ : std_logic;
signal \II_1_counter_13\ : std_logic;
signal \II_1.counter_RNIQ7FB1Z0Z_14\ : std_logic;
signal \II_1_counter_8\ : std_logic;
signal \II_1.counter_RNI6VAM1Z0Z_13_cascade_\ : std_logic;
signal \II_1.counter_RNIJ54VZ0Z_7\ : std_logic;
signal \II_1.counter_RNIA1PIZ0Z_1\ : std_logic;
signal \II_1.counter_RNIJS2EZ0Z_2\ : std_logic;
signal \II_1_counter_12\ : std_logic;
signal \II_1.counter_RNI49153Z0Z_8\ : std_logic;
signal \II_1_counter_27\ : std_logic;
signal \II_1.counter_RNICTOG4Z0Z_12_cascade_\ : std_logic;
signal \II_1.un1_counter_0\ : std_logic;
signal \II_1_counter_26\ : std_logic;
signal \II_1.un1_counterlto22_0\ : std_logic;
signal \II_1.un1_counterlto24_0_0\ : std_logic;
signal \II_1_counter_25\ : std_logic;
signal \II_1_counter_24\ : std_logic;
signal \II_1_counter_23\ : std_logic;
signal \II_1.un1_counterlto25\ : std_logic;
signal \II_1.counterZ0Z_20\ : std_logic;
signal \II_1_counter_19\ : std_logic;
signal \II_1.un1_counterlto25_cascade_\ : std_logic;
signal \II_1_counter_18\ : std_logic;
signal \II_1.counter_RNINVA12Z0Z_20\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PACKAGEPIN_wire\ : std_logic;
signal led6_wire : std_logic;
signal lcol1_wire : std_logic;
signal lcol3_wire : std_logic;
signal led1_wire : std_logic;
signal \PLLOUTGLOBAL_wire\ : std_logic;
signal led2_wire : std_logic;
signal lcol4_wire : std_logic;
signal led4_wire : std_logic;
signal \PLLOUTCORE_wire\ : std_logic;
signal lcol2_wire : std_logic;
signal led7_wire : std_logic;
signal led8_wire : std_logic;
signal led3_wire : std_logic;
signal led5_wire : std_logic;
signal \RESET_wire\ : std_logic;
signal \top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \PACKAGEPIN_wire\ <= PACKAGEPIN;
    led6 <= led6_wire;
    lcol1 <= lcol1_wire;
    lcol3 <= lcol3_wire;
    led1 <= led1_wire;
    PLLOUTGLOBAL <= \PLLOUTGLOBAL_wire\;
    led2 <= led2_wire;
    lcol4 <= lcol4_wire;
    led4 <= led4_wire;
    PLLOUTCORE <= \PLLOUTCORE_wire\;
    lcol2 <= lcol2_wire;
    led7 <= led7_wire;
    led8 <= led8_wire;
    led3 <= led3_wire;
    led5 <= led5_wire;
    \RESET_wire\ <= RESET;
    \top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "010",
            DIVF => "0111000",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => \PLLOUTGLOBAL_0\,
            SDI => '0',
            BYPASS => \GNDG0\,
            RESETB => \N__1298\,
            PLLOUTCORE => \PLLOUTCORE_c\,
            LOCK => OPEN,
            SDO => OPEN,
            SCLK => '0',
            LATCHINPUTVALUE => '0',
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__3086\
        );

    \top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__3086\,
            PACKAGEPIN => \PACKAGEPIN_wire\
        );

    \II_3.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3072\,
            DIN => \N__3071\,
            DOUT => \N__3070\,
            PACKAGEPIN => led6_wire
        );

    \II_3.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__3072\,
            PADOUT => \N__3071\,
            PADIN => \N__3070\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__1372\,
            OUTPUTENABLE => \N__2541\,
            DIN0 => OPEN,
            DOUT0 => \N__1373\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1903\
        );

    \lcol1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3063\,
            DIN => \N__3062\,
            DOUT => \N__3061\,
            PACKAGEPIN => lcol1_wire
        );

    \lcol1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3063\,
            PADOUT => \N__3062\,
            PADIN => \N__3061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3054\,
            DIN => \N__3053\,
            DOUT => \N__3052\,
            PACKAGEPIN => lcol3_wire
        );

    \lcol3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3054\,
            PADOUT => \N__3053\,
            PADIN => \N__3052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2534\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led1_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3045\,
            DIN => \N__3044\,
            DOUT => \N__3043\,
            PACKAGEPIN => led1_wire
        );

    \led1_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3045\,
            PADOUT => \N__3044\,
            PADIN => \N__3043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PLLOUTGLOBAL_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3036\,
            DIN => \N__3035\,
            DOUT => \N__3034\,
            PACKAGEPIN => \PLLOUTGLOBAL_wire\
        );

    \PLLOUTGLOBAL_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3036\,
            PADOUT => \N__3035\,
            PADIN => \N__3034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1337\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led2_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3027\,
            DIN => \N__3026\,
            DOUT => \N__3025\,
            PACKAGEPIN => led2_wire
        );

    \led2_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3027\,
            PADOUT => \N__3026\,
            PADIN => \N__3025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3018\,
            DIN => \N__3017\,
            DOUT => \N__3016\,
            PACKAGEPIN => lcol4_wire
        );

    \lcol4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3018\,
            PADOUT => \N__3017\,
            PADIN => \N__3016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led4_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3009\,
            DIN => \N__3008\,
            DOUT => \N__3007\,
            PACKAGEPIN => led4_wire
        );

    \led4_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3009\,
            PADOUT => \N__3008\,
            PADIN => \N__3007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PLLOUTCORE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3000\,
            DIN => \N__2999\,
            DOUT => \N__2998\,
            PACKAGEPIN => \PLLOUTCORE_wire\
        );

    \PLLOUTCORE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3000\,
            PADOUT => \N__2999\,
            PADIN => \N__2998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1280\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2991\,
            DIN => \N__2990\,
            DOUT => \N__2989\,
            PACKAGEPIN => lcol2_wire
        );

    \lcol2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2991\,
            PADOUT => \N__2990\,
            PADIN => \N__2989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2499\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \II_2.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2982\,
            DIN => \N__2981\,
            DOUT => \N__2980\,
            PACKAGEPIN => led7_wire
        );

    \II_2.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__2982\,
            PADOUT => \N__2981\,
            PADIN => \N__2980\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__1325\,
            OUTPUTENABLE => \N__2558\,
            DIN0 => OPEN,
            DOUT0 => \N__1427\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__1918\
        );

    \led8_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2973\,
            DIN => \N__2972\,
            DOUT => \N__2971\,
            PACKAGEPIN => led8_wire
        );

    \led8_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2973\,
            PADOUT => \N__2972\,
            PADIN => \N__2971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1922\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led3_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2964\,
            DIN => \N__2963\,
            DOUT => \N__2962\,
            PACKAGEPIN => led3_wire
        );

    \led3_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__2964\,
            PADOUT => \N__2963\,
            PADIN => \N__2962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led5_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2955\,
            DIN => \N__2954\,
            DOUT => \N__2953\,
            PACKAGEPIN => led5_wire
        );

    \led5_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__2955\,
            PADOUT => \N__2954\,
            PADIN => \N__2953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESET_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2946\,
            DIN => \N__2945\,
            DOUT => \N__2944\,
            PACKAGEPIN => \RESET_wire\
        );

    \RESET_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2946\,
            PADOUT => \N__2945\,
            PADIN => \N__2944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESET_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__665\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__2924\,
            I => \II_1.counter_RNIA1PIZ0Z_1\
        );

    \I__663\ : InMux
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__661\ : Odrv12
    port map (
            O => \N__2915\,
            I => \II_1.counter_RNIJS2EZ0Z_2\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__659\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2902\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__2908\,
            I => \N__2898\
        );

    \I__657\ : InMux
    port map (
            O => \N__2907\,
            I => \N__2895\
        );

    \I__656\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2892\
        );

    \I__655\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2889\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__2902\,
            I => \N__2886\
        );

    \I__653\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2883\
        );

    \I__652\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2880\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__2895\,
            I => \II_1_counter_12\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__2892\,
            I => \II_1_counter_12\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__2889\,
            I => \II_1_counter_12\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__2886\,
            I => \II_1_counter_12\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__2883\,
            I => \II_1_counter_12\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__2880\,
            I => \II_1_counter_12\
        );

    \I__645\ : InMux
    port map (
            O => \N__2867\,
            I => \N__2864\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__2864\,
            I => \II_1.counter_RNI49153Z0Z_8\
        );

    \I__643\ : InMux
    port map (
            O => \N__2861\,
            I => \N__2857\
        );

    \I__642\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2852\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__2857\,
            I => \N__2849\
        );

    \I__640\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2846\
        );

    \I__639\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2843\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__2852\,
            I => \II_1_counter_27\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__2849\,
            I => \II_1_counter_27\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__2846\,
            I => \II_1_counter_27\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__2843\,
            I => \II_1_counter_27\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__2834\,
            I => \II_1.counter_RNICTOG4Z0Z_12_cascade_\
        );

    \I__633\ : IoInMux
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__2828\,
            I => \II_1.un1_counter_0\
        );

    \I__631\ : InMux
    port map (
            O => \N__2825\,
            I => \N__2821\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__2824\,
            I => \N__2815\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__2821\,
            I => \N__2812\
        );

    \I__628\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2809\
        );

    \I__627\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2804\
        );

    \I__626\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2804\
        );

    \I__625\ : InMux
    port map (
            O => \N__2815\,
            I => \N__2801\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__2812\,
            I => \II_1_counter_26\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__2809\,
            I => \II_1_counter_26\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__2804\,
            I => \II_1_counter_26\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__2801\,
            I => \II_1_counter_26\
        );

    \I__620\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__2789\,
            I => \II_1.un1_counterlto22_0\
        );

    \I__618\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__2783\,
            I => \II_1.un1_counterlto24_0_0\
        );

    \I__616\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2774\
        );

    \I__615\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2771\
        );

    \I__614\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2766\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__2777\,
            I => \N__2762\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2774\,
            I => \N__2757\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__2771\,
            I => \N__2757\
        );

    \I__610\ : InMux
    port map (
            O => \N__2770\,
            I => \N__2754\
        );

    \I__609\ : InMux
    port map (
            O => \N__2769\,
            I => \N__2751\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__2766\,
            I => \N__2748\
        );

    \I__607\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2745\
        );

    \I__606\ : InMux
    port map (
            O => \N__2762\,
            I => \N__2742\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__2757\,
            I => \N__2737\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__2754\,
            I => \N__2737\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__2751\,
            I => \II_1_counter_25\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__2748\,
            I => \II_1_counter_25\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__2745\,
            I => \II_1_counter_25\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__2742\,
            I => \II_1_counter_25\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__2737\,
            I => \II_1_counter_25\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__597\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2719\
        );

    \I__596\ : InMux
    port map (
            O => \N__2722\,
            I => \N__2711\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__2719\,
            I => \N__2708\
        );

    \I__594\ : InMux
    port map (
            O => \N__2718\,
            I => \N__2703\
        );

    \I__593\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2703\
        );

    \I__592\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2700\
        );

    \I__591\ : InMux
    port map (
            O => \N__2715\,
            I => \N__2695\
        );

    \I__590\ : InMux
    port map (
            O => \N__2714\,
            I => \N__2695\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__2711\,
            I => \II_1_counter_24\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__2708\,
            I => \II_1_counter_24\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__2703\,
            I => \II_1_counter_24\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__2700\,
            I => \II_1_counter_24\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__2695\,
            I => \II_1_counter_24\
        );

    \I__584\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2676\
        );

    \I__583\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2673\
        );

    \I__582\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2670\
        );

    \I__581\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2665\
        );

    \I__580\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2665\
        );

    \I__579\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2662\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__2676\,
            I => \II_1_counter_23\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__2673\,
            I => \II_1_counter_23\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__2670\,
            I => \II_1_counter_23\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__2665\,
            I => \II_1_counter_23\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2662\,
            I => \II_1_counter_23\
        );

    \I__573\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2648\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__2648\,
            I => \II_1.un1_counterlto25\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__2645\,
            I => \N__2640\
        );

    \I__570\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2637\
        );

    \I__569\ : InMux
    port map (
            O => \N__2643\,
            I => \N__2634\
        );

    \I__568\ : InMux
    port map (
            O => \N__2640\,
            I => \N__2631\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__2637\,
            I => \N__2628\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__2634\,
            I => \II_1.counterZ0Z_20\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__2631\,
            I => \II_1.counterZ0Z_20\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__2628\,
            I => \II_1.counterZ0Z_20\
        );

    \I__563\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2614\
        );

    \I__562\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2611\
        );

    \I__561\ : InMux
    port map (
            O => \N__2619\,
            I => \N__2606\
        );

    \I__560\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2606\
        );

    \I__559\ : InMux
    port map (
            O => \N__2617\,
            I => \N__2603\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__2614\,
            I => \II_1_counter_19\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__2611\,
            I => \II_1_counter_19\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__2606\,
            I => \II_1_counter_19\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__2603\,
            I => \II_1_counter_19\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__2594\,
            I => \II_1.un1_counterlto25_cascade_\
        );

    \I__553\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2584\
        );

    \I__552\ : InMux
    port map (
            O => \N__2590\,
            I => \N__2581\
        );

    \I__551\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2576\
        );

    \I__550\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2576\
        );

    \I__549\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2573\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2584\,
            I => \II_1_counter_18\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__2581\,
            I => \II_1_counter_18\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2576\,
            I => \II_1_counter_18\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__2573\,
            I => \II_1_counter_18\
        );

    \I__544\ : InMux
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2561\,
            I => \II_1.counter_RNINVA12Z0Z_20\
        );

    \I__542\ : IoInMux
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2555\,
            I => \N__2552\
        );

    \I__540\ : IoSpan4Mux
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__539\ : Span4Mux_s1_v
    port map (
            O => \N__2549\,
            I => \N__2545\
        );

    \I__538\ : IoInMux
    port map (
            O => \N__2548\,
            I => \N__2542\
        );

    \I__537\ : Span4Mux_h
    port map (
            O => \N__2545\,
            I => \N__2535\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2542\,
            I => \N__2535\
        );

    \I__535\ : IoInMux
    port map (
            O => \N__2541\,
            I => \N__2531\
        );

    \I__534\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2528\
        );

    \I__533\ : Span4Mux_s1_v
    port map (
            O => \N__2535\,
            I => \N__2525\
        );

    \I__532\ : IoInMux
    port map (
            O => \N__2534\,
            I => \N__2522\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__2531\,
            I => \N__2519\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__2528\,
            I => \N__2516\
        );

    \I__529\ : Span4Mux_h
    port map (
            O => \N__2525\,
            I => \N__2513\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__2522\,
            I => \N__2510\
        );

    \I__527\ : Span4Mux_s1_v
    port map (
            O => \N__2519\,
            I => \N__2505\
        );

    \I__526\ : Span4Mux_v
    port map (
            O => \N__2516\,
            I => \N__2505\
        );

    \I__525\ : Span4Mux_h
    port map (
            O => \N__2513\,
            I => \N__2500\
        );

    \I__524\ : Span4Mux_s1_v
    port map (
            O => \N__2510\,
            I => \N__2500\
        );

    \I__523\ : Sp12to4
    port map (
            O => \N__2505\,
            I => \N__2494\
        );

    \I__522\ : Sp12to4
    port map (
            O => \N__2500\,
            I => \N__2494\
        );

    \I__521\ : IoInMux
    port map (
            O => \N__2499\,
            I => \N__2491\
        );

    \I__520\ : Span12Mux_h
    port map (
            O => \N__2494\,
            I => \N__2488\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2491\,
            I => \N__2485\
        );

    \I__518\ : Odrv12
    port map (
            O => \N__2488\,
            I => \CONSTANT_ONE_NET\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__2485\,
            I => \CONSTANT_ONE_NET\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__2480\,
            I => \II_3.outputs_RNO_10Z0Z_0_cascade_\
        );

    \I__515\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2474\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2474\,
            I => \N__2471\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__2471\,
            I => \II_3.G_30_0_a3_2_3\
        );

    \I__512\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2463\
        );

    \I__511\ : InMux
    port map (
            O => \N__2467\,
            I => \N__2460\
        );

    \I__510\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2457\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__2463\,
            I => \II_1.counterZ0Z_10\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2460\,
            I => \II_1.counterZ0Z_10\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2457\,
            I => \II_1.counterZ0Z_10\
        );

    \I__506\ : InMux
    port map (
            O => \N__2450\,
            I => \N__2443\
        );

    \I__505\ : InMux
    port map (
            O => \N__2449\,
            I => \N__2440\
        );

    \I__504\ : InMux
    port map (
            O => \N__2448\,
            I => \N__2435\
        );

    \I__503\ : InMux
    port map (
            O => \N__2447\,
            I => \N__2435\
        );

    \I__502\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2432\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2443\,
            I => \II_1_counter_9\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2440\,
            I => \II_1_counter_9\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2435\,
            I => \II_1_counter_9\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__2432\,
            I => \II_1_counter_9\
        );

    \I__497\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2417\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__2422\,
            I => \N__2413\
        );

    \I__495\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2410\
        );

    \I__494\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2407\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2417\,
            I => \N__2404\
        );

    \I__492\ : InMux
    port map (
            O => \N__2416\,
            I => \N__2401\
        );

    \I__491\ : InMux
    port map (
            O => \N__2413\,
            I => \N__2398\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2410\,
            I => \II_1_counter_11\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2407\,
            I => \II_1_counter_11\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__2404\,
            I => \II_1_counter_11\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2401\,
            I => \II_1_counter_11\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2398\,
            I => \II_1_counter_11\
        );

    \I__485\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2382\
        );

    \I__484\ : InMux
    port map (
            O => \N__2386\,
            I => \N__2379\
        );

    \I__483\ : InMux
    port map (
            O => \N__2385\,
            I => \N__2376\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2382\,
            I => \II_1.counterZ0Z_7\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2379\,
            I => \II_1.counterZ0Z_7\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2376\,
            I => \II_1.counterZ0Z_7\
        );

    \I__479\ : InMux
    port map (
            O => \N__2369\,
            I => \N__2362\
        );

    \I__478\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2357\
        );

    \I__477\ : InMux
    port map (
            O => \N__2367\,
            I => \N__2357\
        );

    \I__476\ : InMux
    port map (
            O => \N__2366\,
            I => \N__2352\
        );

    \I__475\ : InMux
    port map (
            O => \N__2365\,
            I => \N__2352\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2362\,
            I => \II_1_counter_16\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__2357\,
            I => \II_1_counter_16\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2352\,
            I => \II_1_counter_16\
        );

    \I__471\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2338\
        );

    \I__470\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2335\
        );

    \I__469\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2332\
        );

    \I__468\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2327\
        );

    \I__467\ : InMux
    port map (
            O => \N__2341\,
            I => \N__2327\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2338\,
            I => \II_1_counter_15\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2335\,
            I => \II_1_counter_15\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2332\,
            I => \II_1_counter_15\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2327\,
            I => \II_1_counter_15\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__2318\,
            I => \N__2311\
        );

    \I__461\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2308\
        );

    \I__460\ : InMux
    port map (
            O => \N__2316\,
            I => \N__2303\
        );

    \I__459\ : InMux
    port map (
            O => \N__2315\,
            I => \N__2303\
        );

    \I__458\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2298\
        );

    \I__457\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2298\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2308\,
            I => \II_1_counter_17\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2303\,
            I => \II_1_counter_17\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2298\,
            I => \II_1_counter_17\
        );

    \I__453\ : InMux
    port map (
            O => \N__2291\,
            I => \N__2287\
        );

    \I__452\ : InMux
    port map (
            O => \N__2290\,
            I => \N__2281\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2287\,
            I => \N__2278\
        );

    \I__450\ : InMux
    port map (
            O => \N__2286\,
            I => \N__2271\
        );

    \I__449\ : InMux
    port map (
            O => \N__2285\,
            I => \N__2271\
        );

    \I__448\ : InMux
    port map (
            O => \N__2284\,
            I => \N__2271\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2281\,
            I => \II_1_counter_14\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__2278\,
            I => \II_1_counter_14\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2271\,
            I => \II_1_counter_14\
        );

    \I__444\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2261\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2261\,
            I => \N__2257\
        );

    \I__442\ : InMux
    port map (
            O => \N__2260\,
            I => \N__2254\
        );

    \I__441\ : Span4Mux_s2_v
    port map (
            O => \N__2257\,
            I => \N__2251\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2254\,
            I => \II_1.counterZ0Z_4\
        );

    \I__439\ : Odrv4
    port map (
            O => \N__2251\,
            I => \II_1.counterZ0Z_4\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__2246\,
            I => \N__2242\
        );

    \I__437\ : InMux
    port map (
            O => \N__2245\,
            I => \N__2238\
        );

    \I__436\ : InMux
    port map (
            O => \N__2242\,
            I => \N__2235\
        );

    \I__435\ : InMux
    port map (
            O => \N__2241\,
            I => \N__2232\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2238\,
            I => \N__2229\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2235\,
            I => \N__2226\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2232\,
            I => \II_1.counterZ0Z_1\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__2229\,
            I => \II_1.counterZ0Z_1\
        );

    \I__430\ : Odrv4
    port map (
            O => \N__2226\,
            I => \II_1.counterZ0Z_1\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__2219\,
            I => \N__2216\
        );

    \I__428\ : InMux
    port map (
            O => \N__2216\,
            I => \N__2212\
        );

    \I__427\ : InMux
    port map (
            O => \N__2215\,
            I => \N__2209\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2212\,
            I => \N__2206\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2209\,
            I => \II_1.counterZ0Z_5\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__2206\,
            I => \II_1.counterZ0Z_5\
        );

    \I__423\ : InMux
    port map (
            O => \N__2201\,
            I => \N__2195\
        );

    \I__422\ : InMux
    port map (
            O => \N__2200\,
            I => \N__2192\
        );

    \I__421\ : InMux
    port map (
            O => \N__2199\,
            I => \N__2187\
        );

    \I__420\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2187\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2195\,
            I => \N__2184\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2192\,
            I => \N__2181\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2187\,
            I => \II_1.counterZ0Z_0\
        );

    \I__416\ : Odrv4
    port map (
            O => \N__2184\,
            I => \II_1.counterZ0Z_0\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__2181\,
            I => \II_1.counterZ0Z_0\
        );

    \I__414\ : InMux
    port map (
            O => \N__2174\,
            I => \N__2169\
        );

    \I__413\ : InMux
    port map (
            O => \N__2173\,
            I => \N__2166\
        );

    \I__412\ : InMux
    port map (
            O => \N__2172\,
            I => \N__2163\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2169\,
            I => \II_1.counterZ0Z_21\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2166\,
            I => \II_1.counterZ0Z_21\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2163\,
            I => \II_1.counterZ0Z_21\
        );

    \I__408\ : InMux
    port map (
            O => \N__2156\,
            I => \N__2149\
        );

    \I__407\ : InMux
    port map (
            O => \N__2155\,
            I => \N__2144\
        );

    \I__406\ : InMux
    port map (
            O => \N__2154\,
            I => \N__2144\
        );

    \I__405\ : InMux
    port map (
            O => \N__2153\,
            I => \N__2139\
        );

    \I__404\ : InMux
    port map (
            O => \N__2152\,
            I => \N__2139\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2149\,
            I => \II_1_counter_22\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2144\,
            I => \II_1_counter_22\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2139\,
            I => \II_1_counter_22\
        );

    \I__400\ : InMux
    port map (
            O => \N__2132\,
            I => \N__2129\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2129\,
            I => \N__2126\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__2126\,
            I => \II_1.un2_clock_outlto23_0_0_c\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__2123\,
            I => \N__2119\
        );

    \I__396\ : InMux
    port map (
            O => \N__2122\,
            I => \N__2113\
        );

    \I__395\ : InMux
    port map (
            O => \N__2119\,
            I => \N__2110\
        );

    \I__394\ : InMux
    port map (
            O => \N__2118\,
            I => \N__2105\
        );

    \I__393\ : InMux
    port map (
            O => \N__2117\,
            I => \N__2105\
        );

    \I__392\ : InMux
    port map (
            O => \N__2116\,
            I => \N__2102\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2113\,
            I => \II_1_counter_13\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2110\,
            I => \II_1_counter_13\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2105\,
            I => \II_1_counter_13\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2102\,
            I => \II_1_counter_13\
        );

    \I__387\ : InMux
    port map (
            O => \N__2093\,
            I => \N__2090\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2090\,
            I => \II_1.counter_RNIQ7FB1Z0Z_14\
        );

    \I__385\ : InMux
    port map (
            O => \N__2087\,
            I => \N__2080\
        );

    \I__384\ : InMux
    port map (
            O => \N__2086\,
            I => \N__2077\
        );

    \I__383\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2074\
        );

    \I__382\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2069\
        );

    \I__381\ : InMux
    port map (
            O => \N__2083\,
            I => \N__2069\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2080\,
            I => \N__2066\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2077\,
            I => \II_1_counter_8\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2074\,
            I => \II_1_counter_8\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2069\,
            I => \II_1_counter_8\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__2066\,
            I => \II_1_counter_8\
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__2057\,
            I => \II_1.counter_RNI6VAM1Z0Z_13_cascade_\
        );

    \I__374\ : InMux
    port map (
            O => \N__2054\,
            I => \N__2051\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2051\,
            I => \II_1.counter_RNIJ54VZ0Z_7\
        );

    \I__372\ : InMux
    port map (
            O => \N__2048\,
            I => \bfn_15_32_0_\
        );

    \I__371\ : InMux
    port map (
            O => \N__2045\,
            I => \II_1.counter_1_cry_25\
        );

    \I__370\ : InMux
    port map (
            O => \N__2042\,
            I => \II_1.counter_1_cry_26\
        );

    \I__369\ : SRMux
    port map (
            O => \N__2039\,
            I => \N__2024\
        );

    \I__368\ : SRMux
    port map (
            O => \N__2038\,
            I => \N__2024\
        );

    \I__367\ : SRMux
    port map (
            O => \N__2037\,
            I => \N__2024\
        );

    \I__366\ : SRMux
    port map (
            O => \N__2036\,
            I => \N__2024\
        );

    \I__365\ : SRMux
    port map (
            O => \N__2035\,
            I => \N__2024\
        );

    \I__364\ : GlobalMux
    port map (
            O => \N__2024\,
            I => \N__2021\
        );

    \I__363\ : gio2CtrlBuf
    port map (
            O => \N__2021\,
            I => \II_1.un1_counter_0_g\
        );

    \I__362\ : InMux
    port map (
            O => \N__2018\,
            I => \N__2013\
        );

    \I__361\ : InMux
    port map (
            O => \N__2017\,
            I => \N__2010\
        );

    \I__360\ : InMux
    port map (
            O => \N__2016\,
            I => \N__2007\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2013\,
            I => \II_1.counterZ0Z_6\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2010\,
            I => \II_1.counterZ0Z_6\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2007\,
            I => \II_1.counterZ0Z_6\
        );

    \I__356\ : InMux
    port map (
            O => \N__2000\,
            I => \N__1996\
        );

    \I__355\ : InMux
    port map (
            O => \N__1999\,
            I => \N__1993\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__1996\,
            I => \II_1.counterZ0Z_2\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__1993\,
            I => \II_1.counterZ0Z_2\
        );

    \I__352\ : InMux
    port map (
            O => \N__1988\,
            I => \N__1984\
        );

    \I__351\ : InMux
    port map (
            O => \N__1987\,
            I => \N__1981\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__1984\,
            I => \II_1.counterZ0Z_3\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__1981\,
            I => \II_1.counterZ0Z_3\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__1976\,
            I => \II_1.un2_clock_outlto19_1_cascade_\
        );

    \I__347\ : InMux
    port map (
            O => \N__1973\,
            I => \N__1970\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__1970\,
            I => \II_1.un2_clock_outlto19_1\
        );

    \I__345\ : InMux
    port map (
            O => \N__1967\,
            I => \N__1964\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__1964\,
            I => \N__1961\
        );

    \I__343\ : Span4Mux_h
    port map (
            O => \N__1961\,
            I => \N__1958\
        );

    \I__342\ : Odrv4
    port map (
            O => \N__1958\,
            I => \II_1.clock_out_RNOZ0Z_3\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__1955\,
            I => \II_1.un2_clock_outlto23_0_0_d_1_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__1952\,
            I => \N__1949\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__1949\,
            I => \N__1945\
        );

    \I__338\ : InMux
    port map (
            O => \N__1948\,
            I => \N__1942\
        );

    \I__337\ : Span4Mux_h
    port map (
            O => \N__1945\,
            I => \N__1938\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1942\,
            I => \N__1935\
        );

    \I__335\ : InMux
    port map (
            O => \N__1941\,
            I => \N__1932\
        );

    \I__334\ : Odrv4
    port map (
            O => \N__1938\,
            I => \counter_RNIG1JB1_20\
        );

    \I__333\ : Odrv4
    port map (
            O => \N__1935\,
            I => \counter_RNIG1JB1_20\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__1932\,
            I => \counter_RNIG1JB1_20\
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__1925\,
            I => \II_1.un2_clock_outlto23_0_0_d_cascade_\
        );

    \I__330\ : IoInMux
    port map (
            O => \N__1922\,
            I => \N__1919\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__1919\,
            I => \N__1915\
        );

    \I__328\ : ClkMux
    port map (
            O => \N__1918\,
            I => \N__1912\
        );

    \I__327\ : IoSpan4Mux
    port map (
            O => \N__1915\,
            I => \N__1907\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1912\,
            I => \N__1907\
        );

    \I__325\ : IoSpan4Mux
    port map (
            O => \N__1907\,
            I => \N__1904\
        );

    \I__324\ : IoSpan4Mux
    port map (
            O => \N__1904\,
            I => \N__1900\
        );

    \I__323\ : ClkMux
    port map (
            O => \N__1903\,
            I => \N__1897\
        );

    \I__322\ : IoSpan4Mux
    port map (
            O => \N__1900\,
            I => \N__1891\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__1897\,
            I => \N__1891\
        );

    \I__320\ : InMux
    port map (
            O => \N__1896\,
            I => \N__1888\
        );

    \I__319\ : IoSpan4Mux
    port map (
            O => \N__1891\,
            I => \N__1885\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1888\,
            I => \N__1882\
        );

    \I__317\ : Span4Mux_s1_v
    port map (
            O => \N__1885\,
            I => \N__1879\
        );

    \I__316\ : Span4Mux_s2_v
    port map (
            O => \N__1882\,
            I => \N__1876\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__1879\,
            I => led8_c
        );

    \I__314\ : Odrv4
    port map (
            O => \N__1876\,
            I => led8_c
        );

    \I__313\ : InMux
    port map (
            O => \N__1871\,
            I => \N__1868\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1868\,
            I => \N__1857\
        );

    \I__311\ : ClkMux
    port map (
            O => \N__1867\,
            I => \N__1838\
        );

    \I__310\ : ClkMux
    port map (
            O => \N__1866\,
            I => \N__1838\
        );

    \I__309\ : ClkMux
    port map (
            O => \N__1865\,
            I => \N__1838\
        );

    \I__308\ : ClkMux
    port map (
            O => \N__1864\,
            I => \N__1838\
        );

    \I__307\ : ClkMux
    port map (
            O => \N__1863\,
            I => \N__1838\
        );

    \I__306\ : ClkMux
    port map (
            O => \N__1862\,
            I => \N__1838\
        );

    \I__305\ : ClkMux
    port map (
            O => \N__1861\,
            I => \N__1838\
        );

    \I__304\ : ClkMux
    port map (
            O => \N__1860\,
            I => \N__1838\
        );

    \I__303\ : Glb2LocalMux
    port map (
            O => \N__1857\,
            I => \N__1838\
        );

    \I__302\ : GlobalMux
    port map (
            O => \N__1838\,
            I => \PLLOUTGLOBAL_0\
        );

    \I__301\ : InMux
    port map (
            O => \N__1835\,
            I => \II_1.counter_1_cry_15\
        );

    \I__300\ : InMux
    port map (
            O => \N__1832\,
            I => \bfn_15_31_0_\
        );

    \I__299\ : InMux
    port map (
            O => \N__1829\,
            I => \II_1.counter_1_cry_17\
        );

    \I__298\ : InMux
    port map (
            O => \N__1826\,
            I => \II_1.counter_1_cry_18\
        );

    \I__297\ : InMux
    port map (
            O => \N__1823\,
            I => \II_1.counter_1_cry_19\
        );

    \I__296\ : InMux
    port map (
            O => \N__1820\,
            I => \II_1.counter_1_cry_20\
        );

    \I__295\ : InMux
    port map (
            O => \N__1817\,
            I => \II_1.counter_1_cry_21\
        );

    \I__294\ : InMux
    port map (
            O => \N__1814\,
            I => \II_1.counter_1_cry_22\
        );

    \I__293\ : InMux
    port map (
            O => \N__1811\,
            I => \II_1.counter_1_cry_23\
        );

    \I__292\ : InMux
    port map (
            O => \N__1808\,
            I => \II_1.counter_1_cry_6\
        );

    \I__291\ : InMux
    port map (
            O => \N__1805\,
            I => \II_1.counter_1_cry_7\
        );

    \I__290\ : InMux
    port map (
            O => \N__1802\,
            I => \bfn_15_30_0_\
        );

    \I__289\ : InMux
    port map (
            O => \N__1799\,
            I => \II_1.counter_1_cry_9\
        );

    \I__288\ : InMux
    port map (
            O => \N__1796\,
            I => \II_1.counter_1_cry_10\
        );

    \I__287\ : InMux
    port map (
            O => \N__1793\,
            I => \II_1.counter_1_cry_11\
        );

    \I__286\ : InMux
    port map (
            O => \N__1790\,
            I => \II_1.counter_1_cry_12\
        );

    \I__285\ : InMux
    port map (
            O => \N__1787\,
            I => \II_1.counter_1_cry_13\
        );

    \I__284\ : InMux
    port map (
            O => \N__1784\,
            I => \II_1.counter_1_cry_14\
        );

    \I__283\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1778\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1778\,
            I => \II_3.G_30_0_o3_0\
        );

    \I__281\ : CascadeMux
    port map (
            O => \N__1775\,
            I => \II_1.counter_RNIM7JB1Z0Z_22_cascade_\
        );

    \I__280\ : InMux
    port map (
            O => \N__1772\,
            I => \N__1769\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1769\,
            I => \N__1766\
        );

    \I__278\ : Odrv4
    port map (
            O => \N__1766\,
            I => \II_1.counter_RNI64GM1Z0Z_26\
        );

    \I__277\ : InMux
    port map (
            O => \N__1763\,
            I => \II_1.counter_1_cry_1\
        );

    \I__276\ : InMux
    port map (
            O => \N__1760\,
            I => \II_1.counter_1_cry_2\
        );

    \I__275\ : InMux
    port map (
            O => \N__1757\,
            I => \II_1.counter_1_cry_3\
        );

    \I__274\ : InMux
    port map (
            O => \N__1754\,
            I => \II_1.counter_1_cry_4\
        );

    \I__273\ : InMux
    port map (
            O => \N__1751\,
            I => \II_1.counter_1_cry_5\
        );

    \I__272\ : InMux
    port map (
            O => \N__1748\,
            I => \N__1745\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1745\,
            I => \II_3.N_14\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__1742\,
            I => \II_3.G_30_0_o3_0_1_cascade_\
        );

    \I__269\ : InMux
    port map (
            O => \N__1739\,
            I => \N__1736\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1736\,
            I => \II_1.counter_RNI1TC9Z0Z_8\
        );

    \I__267\ : InMux
    port map (
            O => \N__1733\,
            I => \N__1730\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1730\,
            I => \II_3.N_16\
        );

    \I__265\ : InMux
    port map (
            O => \N__1727\,
            I => \N__1724\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1724\,
            I => \II_3.G_30_0_a3_1\
        );

    \I__263\ : SRMux
    port map (
            O => \N__1721\,
            I => \N__1718\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1718\,
            I => \N__1715\
        );

    \I__261\ : Odrv4
    port map (
            O => \N__1715\,
            I => \II_3.outputs_RNO_0Z0Z_0\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__1712\,
            I => \N__1706\
        );

    \I__259\ : InMux
    port map (
            O => \N__1711\,
            I => \N__1703\
        );

    \I__258\ : InMux
    port map (
            O => \N__1710\,
            I => \N__1700\
        );

    \I__257\ : InMux
    port map (
            O => \N__1709\,
            I => \N__1695\
        );

    \I__256\ : InMux
    port map (
            O => \N__1706\,
            I => \N__1695\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1703\,
            I => \N__1692\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1700\,
            I => \N__1689\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1695\,
            I => \II_3.counterZ0Z_1\
        );

    \I__252\ : Odrv4
    port map (
            O => \N__1692\,
            I => \II_3.counterZ0Z_1\
        );

    \I__251\ : Odrv4
    port map (
            O => \N__1689\,
            I => \II_3.counterZ0Z_1\
        );

    \I__250\ : CascadeMux
    port map (
            O => \N__1682\,
            I => \N__1678\
        );

    \I__249\ : InMux
    port map (
            O => \N__1681\,
            I => \N__1674\
        );

    \I__248\ : InMux
    port map (
            O => \N__1678\,
            I => \N__1670\
        );

    \I__247\ : InMux
    port map (
            O => \N__1677\,
            I => \N__1667\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1674\,
            I => \N__1664\
        );

    \I__245\ : InMux
    port map (
            O => \N__1673\,
            I => \N__1661\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1670\,
            I => \N__1656\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1667\,
            I => \N__1656\
        );

    \I__242\ : Span4Mux_s1_v
    port map (
            O => \N__1664\,
            I => \N__1653\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1661\,
            I => \II_3.counterZ0Z_2\
        );

    \I__240\ : Odrv4
    port map (
            O => \N__1656\,
            I => \II_3.counterZ0Z_2\
        );

    \I__239\ : Odrv4
    port map (
            O => \N__1653\,
            I => \II_3.counterZ0Z_2\
        );

    \I__238\ : InMux
    port map (
            O => \N__1646\,
            I => \N__1639\
        );

    \I__237\ : InMux
    port map (
            O => \N__1645\,
            I => \N__1636\
        );

    \I__236\ : InMux
    port map (
            O => \N__1644\,
            I => \N__1629\
        );

    \I__235\ : InMux
    port map (
            O => \N__1643\,
            I => \N__1629\
        );

    \I__234\ : InMux
    port map (
            O => \N__1642\,
            I => \N__1629\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1639\,
            I => \N__1626\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1636\,
            I => \N__1623\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1629\,
            I => \II_3.counterZ0Z_0\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__1626\,
            I => \II_3.counterZ0Z_0\
        );

    \I__229\ : Odrv4
    port map (
            O => \N__1623\,
            I => \II_3.counterZ0Z_0\
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__1616\,
            I => \II_3.o2_0_cascade_\
        );

    \I__227\ : CascadeMux
    port map (
            O => \N__1613\,
            I => \N__1610\
        );

    \I__226\ : InMux
    port map (
            O => \N__1610\,
            I => \N__1607\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__1607\,
            I => \II_3.N_12\
        );

    \I__224\ : InMux
    port map (
            O => \N__1604\,
            I => \N__1580\
        );

    \I__223\ : InMux
    port map (
            O => \N__1603\,
            I => \N__1580\
        );

    \I__222\ : InMux
    port map (
            O => \N__1602\,
            I => \N__1580\
        );

    \I__221\ : InMux
    port map (
            O => \N__1601\,
            I => \N__1580\
        );

    \I__220\ : InMux
    port map (
            O => \N__1600\,
            I => \N__1580\
        );

    \I__219\ : InMux
    port map (
            O => \N__1599\,
            I => \N__1580\
        );

    \I__218\ : InMux
    port map (
            O => \N__1598\,
            I => \N__1580\
        );

    \I__217\ : InMux
    port map (
            O => \N__1597\,
            I => \N__1580\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1580\,
            I => \N__1574\
        );

    \I__215\ : InMux
    port map (
            O => \N__1579\,
            I => \N__1571\
        );

    \I__214\ : InMux
    port map (
            O => \N__1578\,
            I => \N__1568\
        );

    \I__213\ : InMux
    port map (
            O => \N__1577\,
            I => \N__1565\
        );

    \I__212\ : Odrv4
    port map (
            O => \N__1574\,
            I => \II_2_G_3_out\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1571\,
            I => \II_2_G_3_out\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1568\,
            I => \II_2_G_3_out\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1565\,
            I => \II_2_G_3_out\
        );

    \I__208\ : CascadeMux
    port map (
            O => \N__1556\,
            I => \N__1550\
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__1555\,
            I => \N__1547\
        );

    \I__206\ : CascadeMux
    port map (
            O => \N__1554\,
            I => \N__1544\
        );

    \I__205\ : InMux
    port map (
            O => \N__1553\,
            I => \N__1533\
        );

    \I__204\ : InMux
    port map (
            O => \N__1550\,
            I => \N__1533\
        );

    \I__203\ : InMux
    port map (
            O => \N__1547\,
            I => \N__1533\
        );

    \I__202\ : InMux
    port map (
            O => \N__1544\,
            I => \N__1533\
        );

    \I__201\ : InMux
    port map (
            O => \N__1543\,
            I => \N__1530\
        );

    \I__200\ : InMux
    port map (
            O => \N__1542\,
            I => \N__1527\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1533\,
            I => \II_2.counterZ0Z_2\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1530\,
            I => \II_2.counterZ0Z_2\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1527\,
            I => \II_2.counterZ0Z_2\
        );

    \I__196\ : CascadeMux
    port map (
            O => \N__1520\,
            I => \N__1516\
        );

    \I__195\ : InMux
    port map (
            O => \N__1519\,
            I => \N__1506\
        );

    \I__194\ : InMux
    port map (
            O => \N__1516\,
            I => \N__1506\
        );

    \I__193\ : InMux
    port map (
            O => \N__1515\,
            I => \N__1506\
        );

    \I__192\ : InMux
    port map (
            O => \N__1514\,
            I => \N__1503\
        );

    \I__191\ : InMux
    port map (
            O => \N__1513\,
            I => \N__1500\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1506\,
            I => \II_2.counterZ0Z_0\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1503\,
            I => \II_2.counterZ0Z_0\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1500\,
            I => \II_2.counterZ0Z_0\
        );

    \I__187\ : InMux
    port map (
            O => \N__1493\,
            I => \N__1482\
        );

    \I__186\ : InMux
    port map (
            O => \N__1492\,
            I => \N__1482\
        );

    \I__185\ : InMux
    port map (
            O => \N__1491\,
            I => \N__1482\
        );

    \I__184\ : InMux
    port map (
            O => \N__1490\,
            I => \N__1479\
        );

    \I__183\ : InMux
    port map (
            O => \N__1489\,
            I => \N__1476\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1482\,
            I => \II_2.counterZ0Z_1\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1479\,
            I => \II_2.counterZ0Z_1\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1476\,
            I => \II_2.counterZ0Z_1\
        );

    \I__179\ : InMux
    port map (
            O => \N__1469\,
            I => \N__1466\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1466\,
            I => \II_2.un1_counter19_1_0\
        );

    \I__177\ : CascadeMux
    port map (
            O => \N__1463\,
            I => \counter_RNI6D8K_6_cascade_\
        );

    \I__176\ : InMux
    port map (
            O => \N__1460\,
            I => \N__1456\
        );

    \I__175\ : InMux
    port map (
            O => \N__1459\,
            I => \N__1453\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1456\,
            I => \counter_RNI6D8K_6\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1453\,
            I => \counter_RNI6D8K_6\
        );

    \I__172\ : CascadeMux
    port map (
            O => \N__1448\,
            I => \II_1.clock_out_RNOZ0Z_5_cascade_\
        );

    \I__171\ : InMux
    port map (
            O => \N__1445\,
            I => \N__1442\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1442\,
            I => \II_1.counter_RNIK1FB1Z0Z_13\
        );

    \I__169\ : InMux
    port map (
            O => \N__1439\,
            I => \N__1436\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1436\,
            I => \II_1.counter_RNIJLJ01_0Z0Z_17\
        );

    \I__167\ : InMux
    port map (
            O => \N__1433\,
            I => \N__1430\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1430\,
            I => \II_1.un1_counterlt12_2\
        );

    \I__165\ : IoInMux
    port map (
            O => \N__1427\,
            I => \N__1424\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1424\,
            I => \N__1421\
        );

    \I__163\ : Span4Mux_s0_v
    port map (
            O => \N__1421\,
            I => \N__1418\
        );

    \I__162\ : Span4Mux_h
    port map (
            O => \N__1418\,
            I => \N__1415\
        );

    \I__161\ : Span4Mux_h
    port map (
            O => \N__1415\,
            I => \N__1411\
        );

    \I__160\ : InMux
    port map (
            O => \N__1414\,
            I => \N__1408\
        );

    \I__159\ : Odrv4
    port map (
            O => \N__1411\,
            I => \II_2.outputsZ0Z_0\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1408\,
            I => \II_2.outputsZ0Z_0\
        );

    \I__157\ : CascadeMux
    port map (
            O => \N__1403\,
            I => \II_1.g3_3_cascade_\
        );

    \I__156\ : CascadeMux
    port map (
            O => \N__1400\,
            I => \II_1.counter_RNIIPRU2Z0Z_11_cascade_\
        );

    \I__155\ : InMux
    port map (
            O => \N__1397\,
            I => \N__1394\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1394\,
            I => \II_1.g0_1_a4_0_0\
        );

    \I__153\ : CEMux
    port map (
            O => \N__1391\,
            I => \N__1388\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1388\,
            I => \N__1385\
        );

    \I__151\ : Span4Mux_v
    port map (
            O => \N__1385\,
            I => \N__1381\
        );

    \I__150\ : InMux
    port map (
            O => \N__1384\,
            I => \N__1378\
        );

    \I__149\ : Odrv4
    port map (
            O => \N__1381\,
            I => \II_1_un2_clock_outlt27_0_i\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1378\,
            I => \II_1_un2_clock_outlt27_0_i\
        );

    \I__147\ : IoInMux
    port map (
            O => \N__1373\,
            I => \N__1369\
        );

    \I__146\ : IoInMux
    port map (
            O => \N__1372\,
            I => \N__1366\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1369\,
            I => \N__1360\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1366\,
            I => \N__1360\
        );

    \I__143\ : InMux
    port map (
            O => \N__1365\,
            I => \N__1357\
        );

    \I__142\ : Odrv4
    port map (
            O => \N__1360\,
            I => \II_3.outputsZ0Z_0\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1357\,
            I => \II_3.outputsZ0Z_0\
        );

    \I__140\ : CascadeMux
    port map (
            O => \N__1352\,
            I => \II_3.o2_cascade_\
        );

    \I__139\ : InMux
    port map (
            O => \N__1349\,
            I => \N__1345\
        );

    \I__138\ : InMux
    port map (
            O => \N__1348\,
            I => \N__1342\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__1345\,
            I => \II_2.un1_counter23_1_5\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__1342\,
            I => \II_2.un1_counter23_1_5\
        );

    \I__135\ : IoInMux
    port map (
            O => \N__1337\,
            I => \N__1334\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__1334\,
            I => \N__1331\
        );

    \I__133\ : Span12Mux_s8_h
    port map (
            O => \N__1331\,
            I => \N__1328\
        );

    \I__132\ : Odrv12
    port map (
            O => \N__1328\,
            I => \GB_BUFFER_PLLOUTGLOBAL_0_THRU_CO\
        );

    \I__131\ : IoInMux
    port map (
            O => \N__1325\,
            I => \N__1322\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__1322\,
            I => \N__1319\
        );

    \I__129\ : IoSpan4Mux
    port map (
            O => \N__1319\,
            I => \N__1316\
        );

    \I__128\ : Span4Mux_s0_v
    port map (
            O => \N__1316\,
            I => \N__1312\
        );

    \I__127\ : CascadeMux
    port map (
            O => \N__1315\,
            I => \N__1309\
        );

    \I__126\ : Span4Mux_h
    port map (
            O => \N__1312\,
            I => \N__1306\
        );

    \I__125\ : InMux
    port map (
            O => \N__1309\,
            I => \N__1303\
        );

    \I__124\ : Odrv4
    port map (
            O => \N__1306\,
            I => \II_2.outputsZ0Z_1\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1303\,
            I => \II_2.outputsZ0Z_1\
        );

    \I__122\ : IoInMux
    port map (
            O => \N__1298\,
            I => \N__1295\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__1295\,
            I => \N__1292\
        );

    \I__120\ : Span12Mux_s7_v
    port map (
            O => \N__1292\,
            I => \N__1289\
        );

    \I__119\ : Span12Mux_h
    port map (
            O => \N__1289\,
            I => \N__1286\
        );

    \I__118\ : Span12Mux_v
    port map (
            O => \N__1286\,
            I => \N__1283\
        );

    \I__117\ : Odrv12
    port map (
            O => \N__1283\,
            I => \RESET_c\
        );

    \I__116\ : IoInMux
    port map (
            O => \N__1280\,
            I => \N__1277\
        );

    \I__115\ : LocalMux
    port map (
            O => \N__1277\,
            I => \N__1274\
        );

    \I__114\ : IoSpan4Mux
    port map (
            O => \N__1274\,
            I => \N__1271\
        );

    \I__113\ : Span4Mux_s3_h
    port map (
            O => \N__1271\,
            I => \N__1268\
        );

    \I__112\ : Sp12to4
    port map (
            O => \N__1268\,
            I => \N__1265\
        );

    \I__111\ : Span12Mux_v
    port map (
            O => \N__1265\,
            I => \N__1262\
        );

    \I__110\ : Span12Mux_h
    port map (
            O => \N__1262\,
            I => \N__1259\
        );

    \I__109\ : Odrv12
    port map (
            O => \N__1259\,
            I => \PLLOUTCORE_c\
        );

    \IN_MUX_bfv_15_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_29_0_\
        );

    \IN_MUX_bfv_15_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \II_1.counter_1_cry_8\,
            carryinitout => \bfn_15_30_0_\
        );

    \IN_MUX_bfv_15_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \II_1.counter_1_cry_16\,
            carryinitout => \bfn_15_31_0_\
        );

    \IN_MUX_bfv_15_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \II_1.counter_1_cry_24\,
            carryinitout => \bfn_15_32_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \II_1.counter_RNIJGA99_0_27\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2831\,
            GLOBALBUFFEROUTPUT => \II_1.un1_counter_0_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \GB_BUFFER_PLLOUTGLOBAL_0_THRU_LUT4_0_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_PLLOUTGLOBAL_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_2.counter_1_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101011110100000"
        )
    port map (
            in0 => \N__1598\,
            in1 => \N__1553\,
            in2 => \N__1520\,
            in3 => \N__1492\,
            lcout => \II_2.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_2.counter_0_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001001111001100"
        )
    port map (
            in0 => \N__1491\,
            in1 => \N__1515\,
            in2 => \N__1555\,
            in3 => \N__1597\,
            lcout => \II_2.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_2.outputs_1_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011110010"
        )
    port map (
            in0 => \N__1601\,
            in1 => \N__1349\,
            in2 => \N__1315\,
            in3 => \N__1469\,
            lcout => \II_2.outputsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_2.counter_2_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__1493\,
            in1 => \N__1519\,
            in2 => \N__1556\,
            in3 => \N__1599\,
            lcout => \II_2.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_3.counter_1_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__1603\,
            in1 => \N__1643\,
            in2 => \_gnd_net_\,
            in3 => \N__1709\,
            lcout => \II_3.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_3.counter_2_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__1644\,
            in1 => \N__1673\,
            in2 => \N__1712\,
            in3 => \N__1604\,
            lcout => \II_3.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_3.counter_0_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__1602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1642\,
            lcout => \II_3.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_2.outputs_0_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110101010"
        )
    port map (
            in0 => \N__1414\,
            in1 => \N__1348\,
            in2 => \N__1554\,
            in3 => \N__1600\,
            lcout => \II_2.outputsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1863\,
            ce => \N__1391\,
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIVSFM1_25_LC_13_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__1941\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2779\,
            lcout => \II_1.g0_1_a4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNI1QAM1_14_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__2540\,
            in1 => \N__1445\,
            in2 => \_gnd_net_\,
            in3 => \N__2291\,
            lcout => OPEN,
            ltout => \II_1.g3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIIPRU2_11_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__1459\,
            in1 => \N__1739\,
            in2 => \N__1403\,
            in3 => \N__2423\,
            lcout => OPEN,
            ltout => \II_1.counter_RNIIPRU2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIAGFC7_11_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100110011"
        )
    port map (
            in0 => \N__1439\,
            in1 => \N__1772\,
            in2 => \N__1400\,
            in3 => \N__1397\,
            lcout => \II_1_un2_clock_outlt27_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_0_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__1365\,
            in1 => \N__1384\,
            in2 => \N__1682\,
            in3 => \N__1579\,
            lcout => \II_3.outputsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1867\,
            ce => 'H',
            sr => \N__1721\
        );

    \II_3.outputs_RNO_5_0_LC_13_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1710\,
            lcout => OPEN,
            ltout => \II_3.o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_1_0_LC_13_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1677\,
            in1 => \N__1645\,
            in2 => \N__1352\,
            in3 => \N__1577\,
            lcout => \II_3.G_30_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_2.counter_RNIEL821_0_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__1542\,
            in1 => \N__1490\,
            in2 => \_gnd_net_\,
            in3 => \N__1514\,
            lcout => \II_2.un1_counter23_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_2.outputs_RNO_0_1_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__1543\,
            in1 => \N__1513\,
            in2 => \_gnd_net_\,
            in3 => \N__1489\,
            lcout => \II_2.un1_counter19_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNI6D8K_6_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2017\,
            in1 => \N__2467\,
            in2 => \_gnd_net_\,
            in3 => \N__2386\,
            lcout => \counter_RNI6D8K_6\,
            ltout => \counter_RNI6D8K_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_9_0_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__2085\,
            in1 => \N__2416\,
            in2 => \N__1463\,
            in3 => \N__2449\,
            lcout => \II_3.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_RNO_5_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2118\,
            in1 => \N__2906\,
            in2 => \_gnd_net_\,
            in3 => \N__2368\,
            lcout => OPEN,
            ltout => \II_1.clock_out_RNOZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_RNO_3_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001111"
        )
    port map (
            in0 => \N__1433\,
            in1 => \N__1460\,
            in2 => \N__1448\,
            in3 => \N__2420\,
            lcout => \II_1.clock_out_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIK1FB1_13_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2117\,
            in1 => \N__2367\,
            in2 => \N__2908\,
            in3 => \N__2343\,
            lcout => \II_1.counter_RNIK1FB1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIJLJ01_0_17_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2619\,
            in1 => \N__2589\,
            in2 => \_gnd_net_\,
            in3 => \N__2316\,
            lcout => \II_1.counter_RNIJLJ01_0Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_RNO_4_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2448\,
            lcout => \II_1.un1_counterlt12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_8_0_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2618\,
            in1 => \N__2588\,
            in2 => \_gnd_net_\,
            in3 => \N__2315\,
            lcout => OPEN,
            ltout => \II_3.G_30_0_o3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_4_0_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__1748\,
            in1 => \N__1948\,
            in2 => \N__1742\,
            in3 => \N__2477\,
            lcout => \II_3.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNI1TC9_8_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2083\,
            lcout => \II_1.counter_RNI1TC9Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_1_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__2199\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2241\,
            lcout => \II_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1865\,
            ce => 'H',
            sr => \N__2037\
        );

    \II_1.counter_RNIG1JB1_20_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__2716\,
            in1 => \N__2682\,
            in2 => \N__2645\,
            in3 => \N__2173\,
            lcout => \counter_RNIG1JB1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_0_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2198\,
            lcout => \II_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1865\,
            ce => 'H',
            sr => \N__2037\
        );

    \II_3.outputs_RNO_0_0_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__1781\,
            in1 => \N__1733\,
            in2 => \N__1613\,
            in3 => \N__1727\,
            lcout => \II_3.outputs_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_6_0_LC_14_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1711\,
            in2 => \_gnd_net_\,
            in3 => \N__2818\,
            lcout => OPEN,
            ltout => \II_3.o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_3_0_LC_14_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1681\,
            in1 => \N__1646\,
            in2 => \N__1616\,
            in3 => \N__1578\,
            lcout => \II_3.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_2.G_3_s_LC_14_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2855\,
            in2 => \_gnd_net_\,
            in3 => \N__1896\,
            lcout => \II_2_G_3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_2_0_LC_14_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__2718\,
            in1 => \N__2681\,
            in2 => \_gnd_net_\,
            in3 => \N__2155\,
            lcout => \II_3.G_30_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIM7JB1_22_LC_14_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__2717\,
            in1 => \N__2680\,
            in2 => \N__2777\,
            in3 => \N__2154\,
            lcout => OPEN,
            ltout => \II_1.counter_RNIM7JB1Z0Z_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNI64GM1_26_LC_14_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1775\,
            in3 => \N__2819\,
            lcout => \II_1.counter_RNI64GM1Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_1_cry_1_c_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2201\,
            in2 => \N__2246\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_29_0_\,
            carryout => \II_1.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_2_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2000\,
            in2 => \_gnd_net_\,
            in3 => \N__1763\,
            lcout => \II_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_1\,
            carryout => \II_1.counter_1_cry_2\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_3_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1988\,
            in2 => \_gnd_net_\,
            in3 => \N__1760\,
            lcout => \II_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_2\,
            carryout => \II_1.counter_1_cry_3\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_4_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2260\,
            in2 => \_gnd_net_\,
            in3 => \N__1757\,
            lcout => \II_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_3\,
            carryout => \II_1.counter_1_cry_4\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_5_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2215\,
            in2 => \_gnd_net_\,
            in3 => \N__1754\,
            lcout => \II_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_4\,
            carryout => \II_1.counter_1_cry_5\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_6_LC_15_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2018\,
            in2 => \_gnd_net_\,
            in3 => \N__1751\,
            lcout => \II_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_5\,
            carryout => \II_1.counter_1_cry_6\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_7_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2387\,
            in2 => \_gnd_net_\,
            in3 => \N__1808\,
            lcout => \II_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_6\,
            carryout => \II_1.counter_1_cry_7\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_8_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2086\,
            in2 => \_gnd_net_\,
            in3 => \N__1805\,
            lcout => \II_1_counter_8\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_7\,
            carryout => \II_1.counter_1_cry_8\,
            clk => \N__1861\,
            ce => 'H',
            sr => \N__2039\
        );

    \II_1.counter_9_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2450\,
            in2 => \_gnd_net_\,
            in3 => \N__1802\,
            lcout => \II_1_counter_9\,
            ltout => OPEN,
            carryin => \bfn_15_30_0_\,
            carryout => \II_1.counter_1_cry_9\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_10_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2468\,
            in2 => \_gnd_net_\,
            in3 => \N__1799\,
            lcout => \II_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_9\,
            carryout => \II_1.counter_1_cry_10\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_11_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2421\,
            in2 => \_gnd_net_\,
            in3 => \N__1796\,
            lcout => \II_1_counter_11\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_10\,
            carryout => \II_1.counter_1_cry_11\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_12_LC_15_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2907\,
            in2 => \_gnd_net_\,
            in3 => \N__1793\,
            lcout => \II_1_counter_12\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_11\,
            carryout => \II_1.counter_1_cry_12\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_13_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2122\,
            in2 => \_gnd_net_\,
            in3 => \N__1790\,
            lcout => \II_1_counter_13\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_12\,
            carryout => \II_1.counter_1_cry_13\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_14_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2290\,
            in2 => \_gnd_net_\,
            in3 => \N__1787\,
            lcout => \II_1_counter_14\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_13\,
            carryout => \II_1.counter_1_cry_14\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_15_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2345\,
            in2 => \_gnd_net_\,
            in3 => \N__1784\,
            lcout => \II_1_counter_15\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_14\,
            carryout => \II_1.counter_1_cry_15\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_16_LC_15_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2369\,
            in2 => \_gnd_net_\,
            in3 => \N__1835\,
            lcout => \II_1_counter_16\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_15\,
            carryout => \II_1.counter_1_cry_16\,
            clk => \N__1862\,
            ce => 'H',
            sr => \N__2038\
        );

    \II_1.counter_17_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2317\,
            in2 => \_gnd_net_\,
            in3 => \N__1832\,
            lcout => \II_1_counter_17\,
            ltout => OPEN,
            carryin => \bfn_15_31_0_\,
            carryout => \II_1.counter_1_cry_17\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_18_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2591\,
            in2 => \_gnd_net_\,
            in3 => \N__1829\,
            lcout => \II_1_counter_18\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_17\,
            carryout => \II_1.counter_1_cry_18\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_19_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2621\,
            in2 => \_gnd_net_\,
            in3 => \N__1826\,
            lcout => \II_1_counter_19\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_18\,
            carryout => \II_1.counter_1_cry_19\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_20_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2643\,
            in2 => \_gnd_net_\,
            in3 => \N__1823\,
            lcout => \II_1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_19\,
            carryout => \II_1.counter_1_cry_20\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_21_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2174\,
            in2 => \_gnd_net_\,
            in3 => \N__1820\,
            lcout => \II_1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_20\,
            carryout => \II_1.counter_1_cry_21\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_22_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2156\,
            in2 => \_gnd_net_\,
            in3 => \N__1817\,
            lcout => \II_1_counter_22\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_21\,
            carryout => \II_1.counter_1_cry_22\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_23_LC_15_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2683\,
            in2 => \_gnd_net_\,
            in3 => \N__1814\,
            lcout => \II_1_counter_23\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_22\,
            carryout => \II_1.counter_1_cry_23\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_24_LC_15_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2722\,
            in2 => \_gnd_net_\,
            in3 => \N__1811\,
            lcout => \II_1_counter_24\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_23\,
            carryout => \II_1.counter_1_cry_24\,
            clk => \N__1864\,
            ce => 'H',
            sr => \N__2036\
        );

    \II_1.counter_25_LC_15_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2769\,
            in2 => \_gnd_net_\,
            in3 => \N__2048\,
            lcout => \II_1_counter_25\,
            ltout => OPEN,
            carryin => \bfn_15_32_0_\,
            carryout => \II_1.counter_1_cry_25\,
            clk => \N__1866\,
            ce => 'H',
            sr => \N__2035\
        );

    \II_1.counter_26_LC_15_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2820\,
            in2 => \_gnd_net_\,
            in3 => \N__2045\,
            lcout => \II_1_counter_26\,
            ltout => OPEN,
            carryin => \II_1.counter_1_cry_25\,
            carryout => \II_1.counter_1_cry_26\,
            clk => \N__1866\,
            ce => 'H',
            sr => \N__2035\
        );

    \II_1.counter_27_LC_15_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2860\,
            in2 => \_gnd_net_\,
            in3 => \N__2042\,
            lcout => \II_1_counter_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1866\,
            ce => 'H',
            sr => \N__2035\
        );

    \II_1.counter_RNIJS2E_2_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2016\,
            in1 => \N__1999\,
            in2 => \_gnd_net_\,
            in3 => \N__1987\,
            lcout => \II_1.counter_RNIJS2EZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIJLJ01_17_LC_16_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2590\,
            in1 => \N__2620\,
            in2 => \_gnd_net_\,
            in3 => \N__2314\,
            lcout => \II_1.un2_clock_outlto19_1\,
            ltout => \II_1.un2_clock_outlto19_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_RNO_2_LC_16_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__2778\,
            in1 => \N__2342\,
            in2 => \N__1976\,
            in3 => \N__2286\,
            lcout => OPEN,
            ltout => \II_1.un2_clock_outlto23_0_0_d_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_RNO_1_LC_16_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111111111"
        )
    port map (
            in0 => \N__1973\,
            in1 => \N__1967\,
            in2 => \N__1955\,
            in3 => \N__1952\,
            lcout => OPEN,
            ltout => \II_1.un2_clock_outlto23_0_0_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_LC_16_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__2132\,
            in1 => \N__2861\,
            in2 => \N__1925\,
            in3 => \N__2825\,
            lcout => led8_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_10_0_LC_16_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2285\,
            in1 => \N__2366\,
            in2 => \N__2123\,
            in3 => \N__2344\,
            lcout => OPEN,
            ltout => \II_3.outputs_RNO_10Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_3.outputs_RNO_7_0_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2480\,
            in3 => \N__2905\,
            lcout => \II_3.G_30_0_a3_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIJ54V_7_LC_16_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2466\,
            in1 => \N__2446\,
            in2 => \N__2422\,
            in3 => \N__2385\,
            lcout => \II_1.counter_RNIJ54VZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIQ7FB1_14_LC_16_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2365\,
            in1 => \N__2341\,
            in2 => \N__2318\,
            in3 => \N__2284\,
            lcout => \II_1.counter_RNIQ7FB1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIA1PI_1_LC_16_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2264\,
            in1 => \N__2245\,
            in2 => \N__2219\,
            in3 => \N__2200\,
            lcout => \II_1.counter_RNIA1PIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNINFPL_21_LC_16_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2152\,
            in2 => \_gnd_net_\,
            in3 => \N__2172\,
            lcout => \II_1.un1_counterlto22_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.clock_out_RNO_0_LC_16_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__2684\,
            in1 => \N__2765\,
            in2 => \N__2726\,
            in3 => \N__2153\,
            lcout => \II_1.un2_clock_outlto23_0_0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNI6VAM1_13_LC_16_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2116\,
            in2 => \_gnd_net_\,
            in3 => \N__2093\,
            lcout => OPEN,
            ltout => \II_1.counter_RNI6VAM1Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNI49153_8_LC_16_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100101"
        )
    port map (
            in0 => \N__2901\,
            in1 => \N__2087\,
            in2 => \N__2057\,
            in3 => \N__2054\,
            lcout => \II_1.counter_RNI49153Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNICTOG4_12_LC_16_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000001111"
        )
    port map (
            in0 => \N__2927\,
            in1 => \N__2921\,
            in2 => \N__2912\,
            in3 => \N__2867\,
            lcout => OPEN,
            ltout => \II_1.counter_RNICTOG4Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIJGA99_27_LC_16_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101010"
        )
    port map (
            in0 => \N__2856\,
            in1 => \N__2564\,
            in2 => \N__2834\,
            in3 => \N__2786\,
            lcout => \II_1.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIVL9C2_26_LC_16_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000011"
        )
    port map (
            in0 => \N__2715\,
            in1 => \N__2651\,
            in2 => \N__2824\,
            in3 => \N__2792\,
            lcout => \II_1.un1_counterlto24_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNIAFM01_23_LC_16_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__2770\,
            in1 => \N__2714\,
            in2 => \_gnd_net_\,
            in3 => \N__2679\,
            lcout => \II_1.un1_counterlto25\,
            ltout => \II_1.un1_counterlto25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \II_1.counter_RNINVA12_20_LC_16_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2644\,
            in1 => \N__2617\,
            in2 => \N__2594\,
            in3 => \N__2587\,
            lcout => \II_1.counter_RNINVA12Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_27_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
