module bum2(PACKAGEPIN,
            PLLOUTCORE,
            PLLOUTGLOBAL,
            RESET);

inout PACKAGEPIN;
input RESET;    /* To initialize the simulation properly, the RESET signal (Active Low) must be asserted at the beginning of the simulation */ 
output PLLOUTCORE;
output PLLOUTGLOBAL;

SB_PLL40_PAD bum2_inst(.PACKAGEPIN(PACKAGEPIN),
                       .PLLOUTCORE(PLLOUTCORE),
                       .PLLOUTGLOBAL(PLLOUTGLOBAL),
                       .EXTFEEDBACK(),
                       .DYNAMICDELAY(),
                       .RESETB(RESET),
                       .BYPASS(1'b0),
                       .LATCHINPUTVALUE(),
                       .LOCK(),
                       .SDI(),
                       .SDO(),
                       .SCLK());

//\\ Fin=12, Fout=171.818;
defparam bum2_inst.DIVR = 4'b0000;
defparam bum2_inst.DIVF = 7'b0111000;
defparam bum2_inst.DIVQ = 3'b010;
defparam bum2_inst.FILTER_RANGE = 3'b001;
defparam bum2_inst.FEEDBACK_PATH = "SIMPLE";
defparam bum2_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
defparam bum2_inst.FDA_FEEDBACK = 4'b0000;
defparam bum2_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
defparam bum2_inst.FDA_RELATIVE = 4'b0000;
defparam bum2_inst.SHIFTREG_DIV_MODE = 2'b00;
defparam bum2_inst.PLLOUT_SELECT = "GENCLK";
defparam bum2_inst.ENABLE_ICEGATE = 1'b0;

endmodule
