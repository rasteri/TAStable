-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 8 2024 23:35:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    led5 : out std_logic;
    lcol2 : out std_logic;
    led6 : out std_logic;
    led2 : out std_logic;
    lcol1 : out std_logic;
    cpuclk : out std_logic;
    apureset : out std_logic;
    led7 : out std_logic;
    led3 : out std_logic;
    lcol4 : out std_logic;
    cpureset : out std_logic;
    apusync : in std_logic;
    PACKAGEPIN : in std_logic;
    masterreset : in std_logic;
    led8 : out std_logic;
    led4 : out std_logic;
    lcol3 : out std_logic;
    led1 : out std_logic;
    consolereset : in std_logic;
    apuclk : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__3600\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2218\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1944\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1902\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1875\ : std_logic;
signal \N__1874\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1840\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1812\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1790\ : std_logic;
signal \N__1787\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1772\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1755\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1728\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1697\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1676\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1641\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1632\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1614\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1586\ : std_logic;
signal \N__1583\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1566\ : std_logic;
signal \N__1563\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1554\ : std_logic;
signal \N__1551\ : std_logic;
signal \N__1548\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1539\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1524\ : std_logic;
signal \N__1521\ : std_logic;
signal \N__1518\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1501\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1498\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1468\ : std_logic;
signal \N__1465\ : std_logic;
signal \N__1462\ : std_logic;
signal \N__1459\ : std_logic;
signal \N__1452\ : std_logic;
signal \N__1443\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1432\ : std_logic;
signal \N__1429\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1423\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1392\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1386\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1380\ : std_logic;
signal \N__1377\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1368\ : std_logic;
signal \top_pll_nrtthrth.PLLOUTCORE_0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \arse.divseven.doutZ0Z_1\ : std_logic;
signal \arse.divseven.N_60_i_cascade_\ : std_logic;
signal \arse.divseven.counter_6_sqmuxa\ : std_logic;
signal \arse.divseven.N_6_cascade_\ : std_logic;
signal \arse.divseven.un1_dout_2_sqmuxa_i_o2_0_cascade_\ : std_logic;
signal \arse.divseven.N_10_cascade_\ : std_logic;
signal \arse.divseven.counterZ0Z_1\ : std_logic;
signal \arse.divseven.counterZ0Z_0\ : std_logic;
signal \arse.divseven.sevenZ0\ : std_logic;
signal \arse.divseven.N_65_i_cascade_\ : std_logic;
signal \arse.divseven.counterZ0Z_2\ : std_logic;
signal \arse.divseven.doutZ0Z_0\ : std_logic;
signal \INVarse.divseven.dout_nesr_0C_net\ : std_logic;
signal \arse.divseven.N_65_i_0\ : std_logic;
signal \arse.seqcounterZ0Z_0\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \arse.seqcounterZ0Z_1\ : std_logic;
signal \arse.un1_seqcounter_1_cry_0\ : std_logic;
signal \arse.seqcounterZ0Z_2\ : std_logic;
signal \arse.un1_seqcounter_1_cry_1\ : std_logic;
signal \arse.seqcounterZ1Z_3\ : std_logic;
signal \arse.un1_seqcounter_1_cry_2\ : std_logic;
signal \arse.un1_seqcounter_1_cry_3\ : std_logic;
signal \arse.seqcounterZ0Z_4\ : std_logic;
signal \arse.seqcounter_i_4\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \arses.un2_counter_cry_1\ : std_logic;
signal \arses.un2_counter_cry_2\ : std_logic;
signal \arses.un2_counter_cry_3\ : std_logic;
signal \arses.counterZ0Z_5\ : std_logic;
signal \arses.un2_counter_cry_4\ : std_logic;
signal \arses.counterZ0Z_6\ : std_logic;
signal \arses.un2_counter_cry_5\ : std_logic;
signal \arses.counterZ0Z_7\ : std_logic;
signal \arses.un2_counter_cry_6\ : std_logic;
signal \arses.counterZ0Z_8\ : std_logic;
signal \arses.un2_counter_cry_7\ : std_logic;
signal \arses.un2_counter_cry_8\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \arses.un2_counter_cry_9\ : std_logic;
signal \arses.un2_counter_cry_10\ : std_logic;
signal \arses.un2_counter_cry_11\ : std_logic;
signal \arses.un2_counter_cry_12\ : std_logic;
signal \arses.un2_counter_cry_13\ : std_logic;
signal \arse.diveight.doutZ0Z_0\ : std_logic;
signal \INVarse.diveight.dout_0C_net\ : std_logic;
signal \arse.diveight.counterZ0Z_1\ : std_logic;
signal \arse.diveight.counterZ0Z_0\ : std_logic;
signal \arses.counterZ0Z_3\ : std_logic;
signal \arses.counterZ0Z_2\ : std_logic;
signal \arses.counterZ0Z_4\ : std_logic;
signal \arses.un1_counterlto4_2_cascade_\ : std_logic;
signal \arses.un1_counterlto8_2\ : std_logic;
signal \arses.counterZ0Z_0\ : std_logic;
signal \arses.counterZ0Z_1\ : std_logic;
signal masterreset_c_i : std_logic;
signal \arses.counterZ0Z_10\ : std_logic;
signal \arses.un1_counterlt11\ : std_logic;
signal \arses.counterZ0Z_11\ : std_logic;
signal \arses.counterZ0Z_9\ : std_logic;
signal \arses.counterZ0Z_14\ : std_logic;
signal \arses.counterZ0Z_13\ : std_logic;
signal \arses.un1_counterlt13_0_cascade_\ : std_logic;
signal \arses.counterZ0Z_12\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \debounceconsolereset.counterZ0Z_2\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_1_THRU_CO\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_1\ : std_logic;
signal \debounceconsolereset.counterZ0Z_3\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_2_THRU_CO\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_2\ : std_logic;
signal \debounceconsolereset.counterZ0Z_4\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_3_THRU_CO\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_3\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_4\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_5\ : std_logic;
signal \clock_out_RNIR6ER_cascade_\ : std_logic;
signal \debounceconsolereset.un1_counterlt6\ : std_logic;
signal masterreset_c : std_logic;
signal \arses.counter8\ : std_logic;
signal \arses.clock_out_i\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_4_THRU_CO\ : std_logic;
signal \debounceconsolereset.counterZ0Z_5\ : std_logic;
signal \debounceconsolereset.out_cnv_3\ : std_logic;
signal \debounceconsolereset.counterZ0Z_6\ : std_logic;
signal consolereset_c : std_logic;
signal \debounceconsolereset.out_cnv_4_cascade_\ : std_logic;
signal \clock_out_RNIR6ER\ : std_logic;
signal \debounceconsolereset.counter_RNI4RTH1Z0Z_6\ : std_logic;
signal \debounceconsolereset.counterZ0Z_0\ : std_logic;
signal \debounceconsolereset.counterZ0Z_1\ : std_logic;
signal \PACKAGEPIN_0_c_g\ : std_logic;
signal \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\ : std_logic;
signal \arse.arse.counterZ0Z_0\ : std_logic;
signal \arse.arse.counterZ0Z_1\ : std_logic;
signal \bfn_16_6_0_\ : std_logic;
signal \arse.arse.counterZ0Z_2\ : std_logic;
signal \arse.arse.un16_counter_cry_1_THRU_CO\ : std_logic;
signal \arse.arse.un16_counter_cry_1\ : std_logic;
signal \arse.arse.un16_counter_cry_2_THRU_CO\ : std_logic;
signal \arse.arse.un16_counter_cry_2\ : std_logic;
signal \arse.arse.un16_counter_cry_3\ : std_logic;
signal \arse.arse.counterZ0Z_4\ : std_logic;
signal \arse.arse.counterZ0Z_3\ : std_logic;
signal \arse.G_2_0_cascade_\ : std_logic;
signal \arse.un1_counterlto4_0\ : std_logic;
signal \arse.un1_counterlt4\ : std_logic;
signal \arse.clock_out_i\ : std_logic;
signal \arse.ddd.Q_esr_RNOZ0Z_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \arse.ddd.N_33_0\ : std_logic;
signal \arse.seqreset_e_0_RNIQTPZ0Z13\ : std_logic;
signal apureset_c : std_logic;
signal \G_73\ : std_logic;
signal apusync_c : std_logic;
signal cpureset_c : std_logic;
signal \arse.seqresetZ0\ : std_logic;
signal \G_74\ : std_logic;
signal \arse.divseven.io_0_D_IN_0\ : std_logic;
signal \G_74_cascade_\ : std_logic;
signal arse_un1_apuclk_i : std_logic;
signal \arse.diveight.counterZ0Z_2\ : std_logic;
signal \arse.diveight.doutZ0Z_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \PLLOUTCORE_0_g\ : std_logic;
signal \arse.seqreset_i\ : std_logic;

signal \PACKAGEPIN_wire\ : std_logic;
signal lcol1_wire : std_logic;
signal masterreset_wire : std_logic;
signal cpureset_wire : std_logic;
signal led8_wire : std_logic;
signal lcol3_wire : std_logic;
signal apuclk_wire : std_logic;
signal lcol4_wire : std_logic;
signal led2_wire : std_logic;
signal led4_wire : std_logic;
signal led6_wire : std_logic;
signal cpuclk_wire : std_logic;
signal apureset_wire : std_logic;
signal consolereset_wire : std_logic;
signal lcol2_wire : std_logic;
signal led1_wire : std_logic;
signal apusync_wire : std_logic;
signal led3_wire : std_logic;
signal led5_wire : std_logic;
signal led7_wire : std_logic;
signal \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \PACKAGEPIN_wire\ <= PACKAGEPIN;
    lcol1 <= lcol1_wire;
    masterreset_wire <= masterreset;
    cpureset <= cpureset_wire;
    led8 <= led8_wire;
    lcol3 <= lcol3_wire;
    apuclk <= apuclk_wire;
    lcol4 <= lcol4_wire;
    led2 <= led2_wire;
    led4 <= led4_wire;
    led6 <= led6_wire;
    cpuclk <= cpuclk_wire;
    apureset <= apureset_wire;
    consolereset_wire <= consolereset;
    lcol2 <= lcol2_wire;
    led1 <= led1_wire;
    apusync_wire <= apusync;
    led3 <= led3_wire;
    led5 <= led5_wire;
    led7 <= led7_wire;
    \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_nrtthrth.top_pll_nrtthrth_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "010",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \top_pll_nrtthrth.PLLOUTCORE_0\,
            REFERENCECLK => \N__2445\,
            RESETB => \N__2318\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PACKAGEPIN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3598\,
            GLOBALBUFFEROUTPUT => \PACKAGEPIN_0_c_g\
        );

    \PACKAGEPIN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3600\,
            DIN => \N__3599\,
            DOUT => \N__3598\,
            PACKAGEPIN => \PACKAGEPIN_wire\
        );

    \PACKAGEPIN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3600\,
            PADOUT => \N__3599\,
            PADIN => \N__3598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3589\,
            DIN => \N__3588\,
            DOUT => \N__3587\,
            PACKAGEPIN => lcol1_wire
        );

    \lcol1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3589\,
            PADOUT => \N__3588\,
            PADIN => \N__3587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \masterreset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3580\,
            DIN => \N__3579\,
            DOUT => \N__3578\,
            PACKAGEPIN => masterreset_wire
        );

    \masterreset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3580\,
            PADOUT => \N__3579\,
            PADIN => \N__3578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => masterreset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \cpureset_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3571\,
            DIN => \N__3570\,
            DOUT => \N__3569\,
            PACKAGEPIN => cpureset_wire
        );

    \cpureset_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3571\,
            PADOUT => \N__3570\,
            PADIN => \N__3569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3177\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3562\,
            DIN => \N__3561\,
            DOUT => \N__3560\,
            PACKAGEPIN => led8_wire
        );

    \led8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3562\,
            PADOUT => \N__3561\,
            PADIN => \N__3560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.divseven.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3553\,
            DIN => \N__3552\,
            DOUT => \N__3551\,
            PACKAGEPIN => OPEN
        );

    \arse.divseven.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__3553\,
            PADOUT => \N__3552\,
            PADIN => \N__3551\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__1398\,
            OUTPUTENABLE => \N__3389\,
            DIN0 => \arse.divseven.io_0_D_IN_0\,
            DOUT0 => \N__1596\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__2933\
        );

    \lcol3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3544\,
            DIN => \N__3543\,
            DOUT => \N__3542\,
            PACKAGEPIN => lcol3_wire
        );

    \lcol3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3544\,
            PADOUT => \N__3543\,
            PADIN => \N__3542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3379\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \apuclk_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3535\,
            DIN => \N__3534\,
            DOUT => \N__3533\,
            PACKAGEPIN => apuclk_wire
        );

    \apuclk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3535\,
            PADOUT => \N__3534\,
            PADIN => \N__3533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3015\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3526\,
            DIN => \N__3525\,
            DOUT => \N__3524\,
            PACKAGEPIN => lcol4_wire
        );

    \lcol4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3526\,
            PADOUT => \N__3525\,
            PADIN => \N__3524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3398\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3517\,
            DIN => \N__3516\,
            DOUT => \N__3515\,
            PACKAGEPIN => led2_wire
        );

    \led2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3517\,
            PADOUT => \N__3516\,
            PADIN => \N__3515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3394\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led4_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3508\,
            DIN => \N__3507\,
            DOUT => \N__3506\,
            PACKAGEPIN => led4_wire
        );

    \led4_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3508\,
            PADOUT => \N__3507\,
            PADIN => \N__3506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led6_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3499\,
            DIN => \N__3498\,
            DOUT => \N__3497\,
            PACKAGEPIN => led6_wire
        );

    \led6_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3499\,
            PADOUT => \N__3498\,
            PADIN => \N__3497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.diveight.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3490\,
            DIN => \N__3489\,
            DOUT => \N__3488\,
            PACKAGEPIN => cpuclk_wire
        );

    \arse.diveight.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__3490\,
            PADOUT => \N__3489\,
            PADIN => \N__3488\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__2958\,
            OUTPUTENABLE => \N__3390\,
            DIN0 => OPEN,
            DOUT0 => \N__1746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__2949\
        );

    \apureset_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3481\,
            DIN => \N__3480\,
            DOUT => \N__3479\,
            PACKAGEPIN => apureset_wire
        );

    \apureset_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3481\,
            PADOUT => \N__3480\,
            PADIN => \N__3479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3268\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \consolereset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3472\,
            DIN => \N__3471\,
            DOUT => \N__3470\,
            PACKAGEPIN => consolereset_wire
        );

    \consolereset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3472\,
            PADOUT => \N__3471\,
            PADIN => \N__3470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => consolereset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3463\,
            DIN => \N__3462\,
            DOUT => \N__3461\,
            PACKAGEPIN => lcol2_wire
        );

    \lcol2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3463\,
            PADOUT => \N__3462\,
            PADIN => \N__3461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3454\,
            DIN => \N__3453\,
            DOUT => \N__3452\,
            PACKAGEPIN => led1_wire
        );

    \led1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3454\,
            PADOUT => \N__3453\,
            PADIN => \N__3452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \apusync_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3445\,
            DIN => \N__3444\,
            DOUT => \N__3443\,
            PACKAGEPIN => apusync_wire
        );

    \apusync_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3445\,
            PADOUT => \N__3444\,
            PADIN => \N__3443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => apusync_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led3_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3436\,
            DIN => \N__3435\,
            DOUT => \N__3434\,
            PACKAGEPIN => led3_wire
        );

    \led3_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3436\,
            PADOUT => \N__3435\,
            PADIN => \N__3434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led5_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3427\,
            DIN => \N__3426\,
            DOUT => \N__3425\,
            PACKAGEPIN => led5_wire
        );

    \led5_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3427\,
            PADOUT => \N__3426\,
            PADIN => \N__3425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led7_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3418\,
            DIN => \N__3417\,
            DOUT => \N__3416\,
            PACKAGEPIN => led7_wire
        );

    \led7_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3418\,
            PADOUT => \N__3417\,
            PADIN => \N__3416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__798\ : IoInMux
    port map (
            O => \N__3399\,
            I => \N__3395\
        );

    \I__797\ : IoInMux
    port map (
            O => \N__3398\,
            I => \N__3391\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__3395\,
            I => \N__3386\
        );

    \I__795\ : IoInMux
    port map (
            O => \N__3394\,
            I => \N__3383\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__3391\,
            I => \N__3380\
        );

    \I__793\ : IoInMux
    port map (
            O => \N__3390\,
            I => \N__3376\
        );

    \I__792\ : IoInMux
    port map (
            O => \N__3389\,
            I => \N__3373\
        );

    \I__791\ : IoSpan4Mux
    port map (
            O => \N__3386\,
            I => \N__3367\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3383\,
            I => \N__3367\
        );

    \I__789\ : IoSpan4Mux
    port map (
            O => \N__3380\,
            I => \N__3364\
        );

    \I__788\ : IoInMux
    port map (
            O => \N__3379\,
            I => \N__3361\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__3376\,
            I => \N__3358\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3355\
        );

    \I__785\ : InMux
    port map (
            O => \N__3372\,
            I => \N__3352\
        );

    \I__784\ : IoSpan4Mux
    port map (
            O => \N__3367\,
            I => \N__3349\
        );

    \I__783\ : IoSpan4Mux
    port map (
            O => \N__3364\,
            I => \N__3344\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__3361\,
            I => \N__3344\
        );

    \I__781\ : IoSpan4Mux
    port map (
            O => \N__3358\,
            I => \N__3341\
        );

    \I__780\ : Span4Mux_s0_h
    port map (
            O => \N__3355\,
            I => \N__3338\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3352\,
            I => \N__3335\
        );

    \I__778\ : IoSpan4Mux
    port map (
            O => \N__3349\,
            I => \N__3330\
        );

    \I__777\ : IoSpan4Mux
    port map (
            O => \N__3344\,
            I => \N__3330\
        );

    \I__776\ : Span4Mux_s3_h
    port map (
            O => \N__3341\,
            I => \N__3327\
        );

    \I__775\ : Span4Mux_h
    port map (
            O => \N__3338\,
            I => \N__3322\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__3335\,
            I => \N__3322\
        );

    \I__773\ : Span4Mux_s2_v
    port map (
            O => \N__3330\,
            I => \N__3319\
        );

    \I__772\ : Sp12to4
    port map (
            O => \N__3327\,
            I => \N__3316\
        );

    \I__771\ : Sp12to4
    port map (
            O => \N__3322\,
            I => \N__3313\
        );

    \I__770\ : Sp12to4
    port map (
            O => \N__3319\,
            I => \N__3310\
        );

    \I__769\ : Span12Mux_h
    port map (
            O => \N__3316\,
            I => \N__3305\
        );

    \I__768\ : Span12Mux_h
    port map (
            O => \N__3313\,
            I => \N__3305\
        );

    \I__767\ : Span12Mux_s8_v
    port map (
            O => \N__3310\,
            I => \N__3302\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__3305\,
            I => \CONSTANT_ONE_NET\
        );

    \I__765\ : Odrv12
    port map (
            O => \N__3302\,
            I => \CONSTANT_ONE_NET\
        );

    \I__764\ : CEMux
    port map (
            O => \N__3297\,
            I => \N__3294\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3294\,
            I => \arse.ddd.N_33_0\
        );

    \I__762\ : SRMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__3285\,
            I => \N__3281\
        );

    \I__759\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3278\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__3281\,
            I => \arse.seqreset_e_0_RNIQTPZ0Z13\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3278\,
            I => \arse.seqreset_e_0_RNIQTPZ0Z13\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__755\ : InMux
    port map (
            O => \N__3270\,
            I => \N__3265\
        );

    \I__754\ : InMux
    port map (
            O => \N__3269\,
            I => \N__3262\
        );

    \I__753\ : IoInMux
    port map (
            O => \N__3268\,
            I => \N__3259\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3265\,
            I => \N__3256\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3262\,
            I => \N__3252\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3259\,
            I => \N__3249\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__3256\,
            I => \N__3246\
        );

    \I__748\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3243\
        );

    \I__747\ : Span4Mux_v
    port map (
            O => \N__3252\,
            I => \N__3240\
        );

    \I__746\ : Span12Mux_s11_h
    port map (
            O => \N__3249\,
            I => \N__3232\
        );

    \I__745\ : Sp12to4
    port map (
            O => \N__3246\,
            I => \N__3232\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3243\,
            I => \N__3232\
        );

    \I__743\ : Span4Mux_h
    port map (
            O => \N__3240\,
            I => \N__3229\
        );

    \I__742\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3226\
        );

    \I__741\ : Odrv12
    port map (
            O => \N__3232\,
            I => apureset_c
        );

    \I__740\ : Odrv4
    port map (
            O => \N__3229\,
            I => apureset_c
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3226\,
            I => apureset_c
        );

    \I__738\ : InMux
    port map (
            O => \N__3219\,
            I => \N__3215\
        );

    \I__737\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3212\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3215\,
            I => \G_73\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3212\,
            I => \G_73\
        );

    \I__734\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3203\
        );

    \I__733\ : InMux
    port map (
            O => \N__3206\,
            I => \N__3200\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3203\,
            I => \N__3194\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3200\,
            I => \N__3194\
        );

    \I__730\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3191\
        );

    \I__729\ : Sp12to4
    port map (
            O => \N__3194\,
            I => \N__3186\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3191\,
            I => \N__3186\
        );

    \I__727\ : Span12Mux_v
    port map (
            O => \N__3186\,
            I => \N__3183\
        );

    \I__726\ : Span12Mux_h
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__3180\,
            I => apusync_c
        );

    \I__724\ : IoInMux
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3174\,
            I => \N__3171\
        );

    \I__722\ : IoSpan4Mux
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__721\ : Span4Mux_s2_h
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__720\ : Span4Mux_h
    port map (
            O => \N__3165\,
            I => \N__3161\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__3164\,
            I => \N__3158\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__3161\,
            I => \N__3155\
        );

    \I__717\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3152\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__3155\,
            I => cpureset_c
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3152\,
            I => cpureset_c
        );

    \I__714\ : InMux
    port map (
            O => \N__3147\,
            I => \N__3143\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__3146\,
            I => \N__3140\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3143\,
            I => \N__3134\
        );

    \I__711\ : InMux
    port map (
            O => \N__3140\,
            I => \N__3131\
        );

    \I__710\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3122\
        );

    \I__709\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3117\
        );

    \I__708\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3117\
        );

    \I__707\ : Span4Mux_v
    port map (
            O => \N__3134\,
            I => \N__3114\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3131\,
            I => \N__3111\
        );

    \I__705\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3108\
        );

    \I__704\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3105\
        );

    \I__703\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3098\
        );

    \I__702\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3098\
        );

    \I__701\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3098\
        );

    \I__700\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3093\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3122\,
            I => \N__3088\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3117\,
            I => \N__3088\
        );

    \I__697\ : Sp12to4
    port map (
            O => \N__3114\,
            I => \N__3083\
        );

    \I__696\ : Span12Mux_s5_v
    port map (
            O => \N__3111\,
            I => \N__3083\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3108\,
            I => \N__3080\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3105\,
            I => \N__3075\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3098\,
            I => \N__3075\
        );

    \I__692\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3069\
        );

    \I__691\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3069\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3093\,
            I => \N__3066\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__3088\,
            I => \N__3063\
        );

    \I__688\ : Span12Mux_h
    port map (
            O => \N__3083\,
            I => \N__3060\
        );

    \I__687\ : Span4Mux_h
    port map (
            O => \N__3080\,
            I => \N__3057\
        );

    \I__686\ : Span12Mux_h
    port map (
            O => \N__3075\,
            I => \N__3054\
        );

    \I__685\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3051\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3069\,
            I => \arse.seqresetZ0\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__3066\,
            I => \arse.seqresetZ0\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__3063\,
            I => \arse.seqresetZ0\
        );

    \I__681\ : Odrv12
    port map (
            O => \N__3060\,
            I => \arse.seqresetZ0\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__3057\,
            I => \arse.seqresetZ0\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__3054\,
            I => \arse.seqresetZ0\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3051\,
            I => \arse.seqresetZ0\
        );

    \I__677\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3033\,
            I => \G_74\
        );

    \I__675\ : InMux
    port map (
            O => \N__3030\,
            I => \N__3027\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3027\,
            I => \N__3024\
        );

    \I__673\ : Span12Mux_h
    port map (
            O => \N__3024\,
            I => \N__3021\
        );

    \I__672\ : Odrv12
    port map (
            O => \N__3021\,
            I => \arse.divseven.io_0_D_IN_0\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__3018\,
            I => \G_74_cascade_\
        );

    \I__670\ : IoInMux
    port map (
            O => \N__3015\,
            I => \N__3012\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3012\,
            I => \N__3009\
        );

    \I__668\ : IoSpan4Mux
    port map (
            O => \N__3009\,
            I => \N__3006\
        );

    \I__667\ : Span4Mux_s3_h
    port map (
            O => \N__3006\,
            I => \N__3003\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__3003\,
            I => \N__3000\
        );

    \I__665\ : Sp12to4
    port map (
            O => \N__3000\,
            I => \N__2997\
        );

    \I__664\ : Odrv12
    port map (
            O => \N__2997\,
            I => arse_un1_apuclk_i
        );

    \I__663\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__2988\,
            I => \N__2985\
        );

    \I__660\ : Sp12to4
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__659\ : Span12Mux_s5_h
    port map (
            O => \N__2982\,
            I => \N__2978\
        );

    \I__658\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2974\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__2978\,
            I => \N__2971\
        );

    \I__656\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2968\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__2974\,
            I => \N__2965\
        );

    \I__654\ : Odrv12
    port map (
            O => \N__2971\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__2968\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__2965\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__651\ : IoInMux
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__2955\,
            I => \N__2952\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__2952\,
            I => \arse.diveight.doutZ0Z_1\
        );

    \I__648\ : ClkMux
    port map (
            O => \N__2949\,
            I => \N__2898\
        );

    \I__647\ : ClkMux
    port map (
            O => \N__2948\,
            I => \N__2898\
        );

    \I__646\ : ClkMux
    port map (
            O => \N__2947\,
            I => \N__2898\
        );

    \I__645\ : ClkMux
    port map (
            O => \N__2946\,
            I => \N__2898\
        );

    \I__644\ : ClkMux
    port map (
            O => \N__2945\,
            I => \N__2898\
        );

    \I__643\ : ClkMux
    port map (
            O => \N__2944\,
            I => \N__2898\
        );

    \I__642\ : ClkMux
    port map (
            O => \N__2943\,
            I => \N__2898\
        );

    \I__641\ : ClkMux
    port map (
            O => \N__2942\,
            I => \N__2898\
        );

    \I__640\ : ClkMux
    port map (
            O => \N__2941\,
            I => \N__2898\
        );

    \I__639\ : ClkMux
    port map (
            O => \N__2940\,
            I => \N__2898\
        );

    \I__638\ : ClkMux
    port map (
            O => \N__2939\,
            I => \N__2898\
        );

    \I__637\ : ClkMux
    port map (
            O => \N__2938\,
            I => \N__2898\
        );

    \I__636\ : ClkMux
    port map (
            O => \N__2937\,
            I => \N__2898\
        );

    \I__635\ : ClkMux
    port map (
            O => \N__2936\,
            I => \N__2898\
        );

    \I__634\ : ClkMux
    port map (
            O => \N__2935\,
            I => \N__2898\
        );

    \I__633\ : ClkMux
    port map (
            O => \N__2934\,
            I => \N__2898\
        );

    \I__632\ : ClkMux
    port map (
            O => \N__2933\,
            I => \N__2898\
        );

    \I__631\ : GlobalMux
    port map (
            O => \N__2898\,
            I => \N__2895\
        );

    \I__630\ : gio2CtrlBuf
    port map (
            O => \N__2895\,
            I => \PLLOUTCORE_0_g\
        );

    \I__629\ : SRMux
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__2889\,
            I => \N__2884\
        );

    \I__627\ : SRMux
    port map (
            O => \N__2888\,
            I => \N__2881\
        );

    \I__626\ : SRMux
    port map (
            O => \N__2887\,
            I => \N__2876\
        );

    \I__625\ : Span4Mux_s3_h
    port map (
            O => \N__2884\,
            I => \N__2873\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__2881\,
            I => \N__2870\
        );

    \I__623\ : SRMux
    port map (
            O => \N__2880\,
            I => \N__2867\
        );

    \I__622\ : SRMux
    port map (
            O => \N__2879\,
            I => \N__2863\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__2876\,
            I => \N__2860\
        );

    \I__620\ : Sp12to4
    port map (
            O => \N__2873\,
            I => \N__2857\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__2870\,
            I => \N__2852\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__2867\,
            I => \N__2852\
        );

    \I__617\ : SRMux
    port map (
            O => \N__2866\,
            I => \N__2849\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__2863\,
            I => \N__2846\
        );

    \I__615\ : Span4Mux_s0_v
    port map (
            O => \N__2860\,
            I => \N__2843\
        );

    \I__614\ : Span12Mux_h
    port map (
            O => \N__2857\,
            I => \N__2834\
        );

    \I__613\ : Sp12to4
    port map (
            O => \N__2852\,
            I => \N__2834\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2849\,
            I => \N__2834\
        );

    \I__611\ : Span4Mux_h
    port map (
            O => \N__2846\,
            I => \N__2831\
        );

    \I__610\ : Span4Mux_h
    port map (
            O => \N__2843\,
            I => \N__2828\
        );

    \I__609\ : SRMux
    port map (
            O => \N__2842\,
            I => \N__2825\
        );

    \I__608\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2822\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__2834\,
            I => \arse.seqreset_i\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__2831\,
            I => \arse.seqreset_i\
        );

    \I__605\ : Odrv4
    port map (
            O => \N__2828\,
            I => \arse.seqreset_i\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__2825\,
            I => \arse.seqreset_i\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__2822\,
            I => \arse.seqreset_i\
        );

    \I__602\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2805\
        );

    \I__601\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2802\
        );

    \I__600\ : InMux
    port map (
            O => \N__2809\,
            I => \N__2799\
        );

    \I__599\ : InMux
    port map (
            O => \N__2808\,
            I => \N__2796\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__2805\,
            I => \arse.arse.counterZ0Z_2\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__2802\,
            I => \arse.arse.counterZ0Z_2\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__2799\,
            I => \arse.arse.counterZ0Z_2\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__2796\,
            I => \arse.arse.counterZ0Z_2\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__2787\,
            I => \N__2784\
        );

    \I__593\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__2781\,
            I => \arse.arse.un16_counter_cry_1_THRU_CO\
        );

    \I__591\ : InMux
    port map (
            O => \N__2778\,
            I => \arse.arse.un16_counter_cry_1\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__2775\,
            I => \N__2772\
        );

    \I__589\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2769\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2769\,
            I => \arse.arse.un16_counter_cry_2_THRU_CO\
        );

    \I__587\ : InMux
    port map (
            O => \N__2766\,
            I => \arse.arse.un16_counter_cry_2\
        );

    \I__586\ : InMux
    port map (
            O => \N__2763\,
            I => \arse.arse.un16_counter_cry_3\
        );

    \I__585\ : InMux
    port map (
            O => \N__2760\,
            I => \N__2756\
        );

    \I__584\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2753\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__2756\,
            I => \arse.arse.counterZ0Z_4\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2753\,
            I => \arse.arse.counterZ0Z_4\
        );

    \I__581\ : InMux
    port map (
            O => \N__2748\,
            I => \N__2743\
        );

    \I__580\ : InMux
    port map (
            O => \N__2747\,
            I => \N__2740\
        );

    \I__579\ : InMux
    port map (
            O => \N__2746\,
            I => \N__2737\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__2743\,
            I => \arse.arse.counterZ0Z_3\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__2740\,
            I => \arse.arse.counterZ0Z_3\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__2737\,
            I => \arse.arse.counterZ0Z_3\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__2730\,
            I => \arse.G_2_0_cascade_\
        );

    \I__574\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2721\
        );

    \I__573\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2721\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__2718\,
            I => \N__2709\
        );

    \I__570\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2706\
        );

    \I__569\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2703\
        );

    \I__568\ : InMux
    port map (
            O => \N__2715\,
            I => \N__2700\
        );

    \I__567\ : InMux
    port map (
            O => \N__2714\,
            I => \N__2693\
        );

    \I__566\ : InMux
    port map (
            O => \N__2713\,
            I => \N__2693\
        );

    \I__565\ : InMux
    port map (
            O => \N__2712\,
            I => \N__2693\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__2709\,
            I => \arse.un1_counterlto4_0\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__2706\,
            I => \arse.un1_counterlto4_0\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__2703\,
            I => \arse.un1_counterlto4_0\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2700\,
            I => \arse.un1_counterlto4_0\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2693\,
            I => \arse.un1_counterlto4_0\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__2682\,
            I => \N__2679\
        );

    \I__558\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2672\
        );

    \I__557\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2663\
        );

    \I__556\ : InMux
    port map (
            O => \N__2677\,
            I => \N__2663\
        );

    \I__555\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2663\
        );

    \I__554\ : InMux
    port map (
            O => \N__2675\,
            I => \N__2660\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__2672\,
            I => \N__2657\
        );

    \I__552\ : InMux
    port map (
            O => \N__2671\,
            I => \N__2652\
        );

    \I__551\ : InMux
    port map (
            O => \N__2670\,
            I => \N__2652\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2663\,
            I => \N__2649\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2660\,
            I => \arse.un1_counterlt4\
        );

    \I__548\ : Odrv4
    port map (
            O => \N__2657\,
            I => \arse.un1_counterlt4\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__2652\,
            I => \arse.un1_counterlt4\
        );

    \I__546\ : Odrv4
    port map (
            O => \N__2649\,
            I => \arse.un1_counterlt4\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__2640\,
            I => \N__2636\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__2639\,
            I => \N__2633\
        );

    \I__543\ : InMux
    port map (
            O => \N__2636\,
            I => \N__2625\
        );

    \I__542\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2625\
        );

    \I__541\ : InMux
    port map (
            O => \N__2632\,
            I => \N__2625\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2625\,
            I => \arse.clock_out_i\
        );

    \I__539\ : InMux
    port map (
            O => \N__2622\,
            I => \N__2619\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__2619\,
            I => \arse.ddd.Q_esr_RNOZ0Z_0\
        );

    \I__537\ : InMux
    port map (
            O => \N__2616\,
            I => \N__2613\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__535\ : Span12Mux_v
    port map (
            O => \N__2610\,
            I => \N__2607\
        );

    \I__534\ : Span12Mux_v
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__533\ : Odrv12
    port map (
            O => \N__2604\,
            I => consolereset_c
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__2601\,
            I => \debounceconsolereset.out_cnv_4_cascade_\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__2598\,
            I => \N__2592\
        );

    \I__530\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2583\
        );

    \I__529\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2583\
        );

    \I__528\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2580\
        );

    \I__527\ : InMux
    port map (
            O => \N__2592\,
            I => \N__2575\
        );

    \I__526\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2575\
        );

    \I__525\ : InMux
    port map (
            O => \N__2590\,
            I => \N__2568\
        );

    \I__524\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2568\
        );

    \I__523\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2568\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2583\,
            I => \clock_out_RNIR6ER\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__2580\,
            I => \clock_out_RNIR6ER\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__2575\,
            I => \clock_out_RNIR6ER\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2568\,
            I => \clock_out_RNIR6ER\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__2559\,
            I => \N__2556\
        );

    \I__517\ : InMux
    port map (
            O => \N__2556\,
            I => \N__2547\
        );

    \I__516\ : InMux
    port map (
            O => \N__2555\,
            I => \N__2542\
        );

    \I__515\ : InMux
    port map (
            O => \N__2554\,
            I => \N__2542\
        );

    \I__514\ : InMux
    port map (
            O => \N__2553\,
            I => \N__2533\
        );

    \I__513\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2533\
        );

    \I__512\ : InMux
    port map (
            O => \N__2551\,
            I => \N__2533\
        );

    \I__511\ : InMux
    port map (
            O => \N__2550\,
            I => \N__2533\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2547\,
            I => \debounceconsolereset.counter_RNI4RTH1Z0Z_6\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__2542\,
            I => \debounceconsolereset.counter_RNI4RTH1Z0Z_6\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2533\,
            I => \debounceconsolereset.counter_RNI4RTH1Z0Z_6\
        );

    \I__507\ : InMux
    port map (
            O => \N__2526\,
            I => \N__2522\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__2525\,
            I => \N__2517\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__2522\,
            I => \N__2514\
        );

    \I__504\ : InMux
    port map (
            O => \N__2521\,
            I => \N__2509\
        );

    \I__503\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2509\
        );

    \I__502\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2506\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__2514\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2509\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2506\,
            I => \debounceconsolereset.counterZ0Z_0\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__2499\,
            I => \N__2495\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__2498\,
            I => \N__2492\
        );

    \I__496\ : InMux
    port map (
            O => \N__2495\,
            I => \N__2486\
        );

    \I__495\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2486\
        );

    \I__494\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2483\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2486\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2483\,
            I => \debounceconsolereset.counterZ0Z_1\
        );

    \I__491\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2475\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2475\,
            I => \N__2466\
        );

    \I__489\ : ClkMux
    port map (
            O => \N__2474\,
            I => \N__2451\
        );

    \I__488\ : ClkMux
    port map (
            O => \N__2473\,
            I => \N__2451\
        );

    \I__487\ : ClkMux
    port map (
            O => \N__2472\,
            I => \N__2451\
        );

    \I__486\ : ClkMux
    port map (
            O => \N__2471\,
            I => \N__2451\
        );

    \I__485\ : ClkMux
    port map (
            O => \N__2470\,
            I => \N__2451\
        );

    \I__484\ : ClkMux
    port map (
            O => \N__2469\,
            I => \N__2451\
        );

    \I__483\ : Glb2LocalMux
    port map (
            O => \N__2466\,
            I => \N__2451\
        );

    \I__482\ : GlobalMux
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__481\ : gio2CtrlBuf
    port map (
            O => \N__2448\,
            I => \PACKAGEPIN_0_c_g\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__2445\,
            I => \N__2442\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2442\,
            I => \N__2439\
        );

    \I__478\ : IoSpan4Mux
    port map (
            O => \N__2439\,
            I => \N__2436\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__2436\,
            I => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\
        );

    \I__476\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2427\
        );

    \I__475\ : InMux
    port map (
            O => \N__2432\,
            I => \N__2424\
        );

    \I__474\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2421\
        );

    \I__473\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2418\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2427\,
            I => \arse.arse.counterZ0Z_0\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2424\,
            I => \arse.arse.counterZ0Z_0\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2421\,
            I => \arse.arse.counterZ0Z_0\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2418\,
            I => \arse.arse.counterZ0Z_0\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2409\,
            I => \N__2405\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__2408\,
            I => \N__2402\
        );

    \I__466\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2398\
        );

    \I__465\ : InMux
    port map (
            O => \N__2402\,
            I => \N__2395\
        );

    \I__464\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2392\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2398\,
            I => \arse.arse.counterZ0Z_1\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2395\,
            I => \arse.arse.counterZ0Z_1\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__2392\,
            I => \arse.arse.counterZ0Z_1\
        );

    \I__460\ : InMux
    port map (
            O => \N__2385\,
            I => \N__2382\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2382\,
            I => \debounceconsolereset.un3_counter_cry_2_THRU_CO\
        );

    \I__458\ : InMux
    port map (
            O => \N__2379\,
            I => \debounceconsolereset.un3_counter_cry_2\
        );

    \I__457\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2370\
        );

    \I__456\ : InMux
    port map (
            O => \N__2375\,
            I => \N__2363\
        );

    \I__455\ : InMux
    port map (
            O => \N__2374\,
            I => \N__2363\
        );

    \I__454\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2363\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2370\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2363\,
            I => \debounceconsolereset.counterZ0Z_4\
        );

    \I__451\ : InMux
    port map (
            O => \N__2358\,
            I => \N__2355\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2355\,
            I => \debounceconsolereset.un3_counter_cry_3_THRU_CO\
        );

    \I__449\ : InMux
    port map (
            O => \N__2352\,
            I => \debounceconsolereset.un3_counter_cry_3\
        );

    \I__448\ : InMux
    port map (
            O => \N__2349\,
            I => \debounceconsolereset.un3_counter_cry_4\
        );

    \I__447\ : InMux
    port map (
            O => \N__2346\,
            I => \debounceconsolereset.un3_counter_cry_5\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__2343\,
            I => \clock_out_RNIR6ER_cascade_\
        );

    \I__445\ : InMux
    port map (
            O => \N__2340\,
            I => \N__2337\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2337\,
            I => \debounceconsolereset.un1_counterlt6\
        );

    \I__443\ : InMux
    port map (
            O => \N__2334\,
            I => \N__2330\
        );

    \I__442\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2327\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2330\,
            I => \N__2322\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2327\,
            I => \N__2319\
        );

    \I__439\ : InMux
    port map (
            O => \N__2326\,
            I => \N__2315\
        );

    \I__438\ : CEMux
    port map (
            O => \N__2325\,
            I => \N__2312\
        );

    \I__437\ : Span4Mux_v
    port map (
            O => \N__2322\,
            I => \N__2304\
        );

    \I__436\ : Span4Mux_v
    port map (
            O => \N__2319\,
            I => \N__2301\
        );

    \I__435\ : IoInMux
    port map (
            O => \N__2318\,
            I => \N__2298\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2315\,
            I => \N__2295\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2312\,
            I => \N__2292\
        );

    \I__432\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2285\
        );

    \I__431\ : InMux
    port map (
            O => \N__2310\,
            I => \N__2285\
        );

    \I__430\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2285\
        );

    \I__429\ : InMux
    port map (
            O => \N__2308\,
            I => \N__2280\
        );

    \I__428\ : InMux
    port map (
            O => \N__2307\,
            I => \N__2280\
        );

    \I__427\ : Span4Mux_h
    port map (
            O => \N__2304\,
            I => \N__2275\
        );

    \I__426\ : Span4Mux_h
    port map (
            O => \N__2301\,
            I => \N__2275\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2298\,
            I => \N__2272\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__2295\,
            I => \N__2269\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__2292\,
            I => \N__2262\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2285\,
            I => \N__2262\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2280\,
            I => \N__2262\
        );

    \I__420\ : Span4Mux_h
    port map (
            O => \N__2275\,
            I => \N__2257\
        );

    \I__419\ : Span4Mux_s2_v
    port map (
            O => \N__2272\,
            I => \N__2257\
        );

    \I__418\ : Sp12to4
    port map (
            O => \N__2269\,
            I => \N__2254\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__2262\,
            I => \N__2251\
        );

    \I__416\ : Span4Mux_h
    port map (
            O => \N__2257\,
            I => \N__2248\
        );

    \I__415\ : Span12Mux_h
    port map (
            O => \N__2254\,
            I => \N__2245\
        );

    \I__414\ : Sp12to4
    port map (
            O => \N__2251\,
            I => \N__2242\
        );

    \I__413\ : Span4Mux_h
    port map (
            O => \N__2248\,
            I => \N__2239\
        );

    \I__412\ : Span12Mux_h
    port map (
            O => \N__2245\,
            I => \N__2236\
        );

    \I__411\ : Span12Mux_h
    port map (
            O => \N__2242\,
            I => \N__2233\
        );

    \I__410\ : Sp12to4
    port map (
            O => \N__2239\,
            I => \N__2230\
        );

    \I__409\ : Span12Mux_v
    port map (
            O => \N__2236\,
            I => \N__2227\
        );

    \I__408\ : Span12Mux_h
    port map (
            O => \N__2233\,
            I => \N__2224\
        );

    \I__407\ : Span12Mux_v
    port map (
            O => \N__2230\,
            I => \N__2221\
        );

    \I__406\ : Span12Mux_v
    port map (
            O => \N__2227\,
            I => \N__2218\
        );

    \I__405\ : Span12Mux_v
    port map (
            O => \N__2224\,
            I => \N__2215\
        );

    \I__404\ : Span12Mux_v
    port map (
            O => \N__2221\,
            I => \N__2212\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__2218\,
            I => masterreset_c
        );

    \I__402\ : Odrv12
    port map (
            O => \N__2215\,
            I => masterreset_c
        );

    \I__401\ : Odrv12
    port map (
            O => \N__2212\,
            I => masterreset_c
        );

    \I__400\ : InMux
    port map (
            O => \N__2205\,
            I => \N__2186\
        );

    \I__399\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2177\
        );

    \I__398\ : InMux
    port map (
            O => \N__2203\,
            I => \N__2177\
        );

    \I__397\ : InMux
    port map (
            O => \N__2202\,
            I => \N__2177\
        );

    \I__396\ : InMux
    port map (
            O => \N__2201\,
            I => \N__2177\
        );

    \I__395\ : InMux
    port map (
            O => \N__2200\,
            I => \N__2170\
        );

    \I__394\ : InMux
    port map (
            O => \N__2199\,
            I => \N__2170\
        );

    \I__393\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2170\
        );

    \I__392\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2165\
        );

    \I__391\ : InMux
    port map (
            O => \N__2196\,
            I => \N__2165\
        );

    \I__390\ : InMux
    port map (
            O => \N__2195\,
            I => \N__2158\
        );

    \I__389\ : InMux
    port map (
            O => \N__2194\,
            I => \N__2158\
        );

    \I__388\ : InMux
    port map (
            O => \N__2193\,
            I => \N__2158\
        );

    \I__387\ : InMux
    port map (
            O => \N__2192\,
            I => \N__2151\
        );

    \I__386\ : InMux
    port map (
            O => \N__2191\,
            I => \N__2151\
        );

    \I__385\ : InMux
    port map (
            O => \N__2190\,
            I => \N__2151\
        );

    \I__384\ : InMux
    port map (
            O => \N__2189\,
            I => \N__2148\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2186\,
            I => \arses.counter8\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2177\,
            I => \arses.counter8\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2170\,
            I => \arses.counter8\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2165\,
            I => \arses.counter8\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2158\,
            I => \arses.counter8\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2151\,
            I => \arses.counter8\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2148\,
            I => \arses.counter8\
        );

    \I__376\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2129\
        );

    \I__375\ : InMux
    port map (
            O => \N__2132\,
            I => \N__2126\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2129\,
            I => \arses.clock_out_i\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2126\,
            I => \arses.clock_out_i\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2121\,
            I => \N__2118\
        );

    \I__371\ : InMux
    port map (
            O => \N__2118\,
            I => \N__2115\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2115\,
            I => \debounceconsolereset.un3_counter_cry_4_THRU_CO\
        );

    \I__369\ : InMux
    port map (
            O => \N__2112\,
            I => \N__2104\
        );

    \I__368\ : InMux
    port map (
            O => \N__2111\,
            I => \N__2104\
        );

    \I__367\ : InMux
    port map (
            O => \N__2110\,
            I => \N__2099\
        );

    \I__366\ : InMux
    port map (
            O => \N__2109\,
            I => \N__2099\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2104\,
            I => \debounceconsolereset.counterZ0Z_5\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2099\,
            I => \debounceconsolereset.counterZ0Z_5\
        );

    \I__363\ : InMux
    port map (
            O => \N__2094\,
            I => \N__2091\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2091\,
            I => \N__2088\
        );

    \I__361\ : Odrv4
    port map (
            O => \N__2088\,
            I => \debounceconsolereset.out_cnv_3\
        );

    \I__360\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2080\
        );

    \I__359\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2077\
        );

    \I__358\ : InMux
    port map (
            O => \N__2083\,
            I => \N__2074\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2080\,
            I => \debounceconsolereset.counterZ0Z_6\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2077\,
            I => \debounceconsolereset.counterZ0Z_6\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2074\,
            I => \debounceconsolereset.counterZ0Z_6\
        );

    \I__354\ : InMux
    port map (
            O => \N__2067\,
            I => \N__2063\
        );

    \I__353\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2060\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2063\,
            I => \arses.counterZ0Z_14\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2060\,
            I => \arses.counterZ0Z_14\
        );

    \I__350\ : InMux
    port map (
            O => \N__2055\,
            I => \N__2051\
        );

    \I__349\ : InMux
    port map (
            O => \N__2054\,
            I => \N__2048\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2051\,
            I => \arses.counterZ0Z_13\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2048\,
            I => \arses.counterZ0Z_13\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__2043\,
            I => \arses.un1_counterlt13_0_cascade_\
        );

    \I__345\ : InMux
    port map (
            O => \N__2040\,
            I => \N__2036\
        );

    \I__344\ : InMux
    port map (
            O => \N__2039\,
            I => \N__2033\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2036\,
            I => \arses.counterZ0Z_12\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2033\,
            I => \arses.counterZ0Z_12\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2028\,
            I => \N__2025\
        );

    \I__340\ : InMux
    port map (
            O => \N__2025\,
            I => \N__2015\
        );

    \I__339\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2015\
        );

    \I__338\ : InMux
    port map (
            O => \N__2023\,
            I => \N__2015\
        );

    \I__337\ : InMux
    port map (
            O => \N__2022\,
            I => \N__2012\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2015\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2012\,
            I => \debounceconsolereset.counterZ0Z_2\
        );

    \I__334\ : InMux
    port map (
            O => \N__2007\,
            I => \N__2004\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2004\,
            I => \debounceconsolereset.un3_counter_cry_1_THRU_CO\
        );

    \I__332\ : InMux
    port map (
            O => \N__2001\,
            I => \debounceconsolereset.un3_counter_cry_1\
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__1998\,
            I => \N__1993\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__1997\,
            I => \N__1990\
        );

    \I__329\ : InMux
    port map (
            O => \N__1996\,
            I => \N__1986\
        );

    \I__328\ : InMux
    port map (
            O => \N__1993\,
            I => \N__1979\
        );

    \I__327\ : InMux
    port map (
            O => \N__1990\,
            I => \N__1979\
        );

    \I__326\ : InMux
    port map (
            O => \N__1989\,
            I => \N__1979\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__1986\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1979\,
            I => \debounceconsolereset.counterZ0Z_3\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__1974\,
            I => \N__1971\
        );

    \I__322\ : InMux
    port map (
            O => \N__1971\,
            I => \N__1965\
        );

    \I__321\ : InMux
    port map (
            O => \N__1970\,
            I => \N__1965\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__1965\,
            I => \arse.diveight.counterZ0Z_1\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__1962\,
            I => \N__1958\
        );

    \I__318\ : InMux
    port map (
            O => \N__1961\,
            I => \N__1954\
        );

    \I__317\ : InMux
    port map (
            O => \N__1958\,
            I => \N__1949\
        );

    \I__316\ : InMux
    port map (
            O => \N__1957\,
            I => \N__1949\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__1954\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__1949\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__313\ : InMux
    port map (
            O => \N__1944\,
            I => \N__1940\
        );

    \I__312\ : InMux
    port map (
            O => \N__1943\,
            I => \N__1937\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__1940\,
            I => \arses.counterZ0Z_3\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1937\,
            I => \arses.counterZ0Z_3\
        );

    \I__309\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1928\
        );

    \I__308\ : InMux
    port map (
            O => \N__1931\,
            I => \N__1925\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1928\,
            I => \arses.counterZ0Z_2\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1925\,
            I => \arses.counterZ0Z_2\
        );

    \I__305\ : InMux
    port map (
            O => \N__1920\,
            I => \N__1916\
        );

    \I__304\ : InMux
    port map (
            O => \N__1919\,
            I => \N__1913\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1916\,
            I => \N__1910\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1913\,
            I => \arses.counterZ0Z_4\
        );

    \I__301\ : Odrv4
    port map (
            O => \N__1910\,
            I => \arses.counterZ0Z_4\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__1905\,
            I => \arses.un1_counterlto4_2_cascade_\
        );

    \I__299\ : InMux
    port map (
            O => \N__1902\,
            I => \N__1899\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1899\,
            I => \arses.un1_counterlto8_2\
        );

    \I__297\ : InMux
    port map (
            O => \N__1896\,
            I => \N__1893\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1893\,
            I => \N__1887\
        );

    \I__295\ : InMux
    port map (
            O => \N__1892\,
            I => \N__1880\
        );

    \I__294\ : InMux
    port map (
            O => \N__1891\,
            I => \N__1880\
        );

    \I__293\ : InMux
    port map (
            O => \N__1890\,
            I => \N__1880\
        );

    \I__292\ : Odrv4
    port map (
            O => \N__1887\,
            I => \arses.counterZ0Z_0\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1880\,
            I => \arses.counterZ0Z_0\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__1875\,
            I => \N__1871\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__1874\,
            I => \N__1868\
        );

    \I__288\ : InMux
    port map (
            O => \N__1871\,
            I => \N__1864\
        );

    \I__287\ : InMux
    port map (
            O => \N__1868\,
            I => \N__1859\
        );

    \I__286\ : InMux
    port map (
            O => \N__1867\,
            I => \N__1859\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1864\,
            I => \arses.counterZ0Z_1\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1859\,
            I => \arses.counterZ0Z_1\
        );

    \I__283\ : SRMux
    port map (
            O => \N__1854\,
            I => \N__1849\
        );

    \I__282\ : SRMux
    port map (
            O => \N__1853\,
            I => \N__1846\
        );

    \I__281\ : SRMux
    port map (
            O => \N__1852\,
            I => \N__1843\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1849\,
            I => \N__1840\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1846\,
            I => \N__1835\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1843\,
            I => \N__1835\
        );

    \I__277\ : Span4Mux_v
    port map (
            O => \N__1840\,
            I => \N__1832\
        );

    \I__276\ : Odrv4
    port map (
            O => \N__1835\,
            I => masterreset_c_i
        );

    \I__275\ : Odrv4
    port map (
            O => \N__1832\,
            I => masterreset_c_i
        );

    \I__274\ : InMux
    port map (
            O => \N__1827\,
            I => \N__1823\
        );

    \I__273\ : InMux
    port map (
            O => \N__1826\,
            I => \N__1820\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1823\,
            I => \arses.counterZ0Z_10\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1820\,
            I => \arses.counterZ0Z_10\
        );

    \I__270\ : InMux
    port map (
            O => \N__1815\,
            I => \N__1812\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1812\,
            I => \arses.un1_counterlt11\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__1809\,
            I => \N__1805\
        );

    \I__267\ : InMux
    port map (
            O => \N__1808\,
            I => \N__1802\
        );

    \I__266\ : InMux
    port map (
            O => \N__1805\,
            I => \N__1799\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1802\,
            I => \arses.counterZ0Z_11\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1799\,
            I => \arses.counterZ0Z_11\
        );

    \I__263\ : InMux
    port map (
            O => \N__1794\,
            I => \N__1790\
        );

    \I__262\ : InMux
    port map (
            O => \N__1793\,
            I => \N__1787\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1790\,
            I => \arses.counterZ0Z_9\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__1787\,
            I => \arses.counterZ0Z_9\
        );

    \I__259\ : CascadeMux
    port map (
            O => \N__1782\,
            I => \N__1778\
        );

    \I__258\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1775\
        );

    \I__257\ : InMux
    port map (
            O => \N__1778\,
            I => \N__1772\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1775\,
            I => \arses.counterZ0Z_8\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1772\,
            I => \arses.counterZ0Z_8\
        );

    \I__254\ : InMux
    port map (
            O => \N__1767\,
            I => \arses.un2_counter_cry_7\
        );

    \I__253\ : InMux
    port map (
            O => \N__1764\,
            I => \bfn_9_5_0_\
        );

    \I__252\ : InMux
    port map (
            O => \N__1761\,
            I => \arses.un2_counter_cry_9\
        );

    \I__251\ : InMux
    port map (
            O => \N__1758\,
            I => \arses.un2_counter_cry_10\
        );

    \I__250\ : InMux
    port map (
            O => \N__1755\,
            I => \arses.un2_counter_cry_11\
        );

    \I__249\ : InMux
    port map (
            O => \N__1752\,
            I => \arses.un2_counter_cry_12\
        );

    \I__248\ : InMux
    port map (
            O => \N__1749\,
            I => \arses.un2_counter_cry_13\
        );

    \I__247\ : IoInMux
    port map (
            O => \N__1746\,
            I => \N__1743\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1743\,
            I => \N__1740\
        );

    \I__245\ : Span4Mux_s1_h
    port map (
            O => \N__1740\,
            I => \N__1737\
        );

    \I__244\ : Span4Mux_v
    port map (
            O => \N__1737\,
            I => \N__1734\
        );

    \I__243\ : Sp12to4
    port map (
            O => \N__1734\,
            I => \N__1731\
        );

    \I__242\ : Span12Mux_h
    port map (
            O => \N__1731\,
            I => \N__1728\
        );

    \I__241\ : Odrv12
    port map (
            O => \N__1728\,
            I => \arse.diveight.doutZ0Z_0\
        );

    \I__240\ : InMux
    port map (
            O => \N__1725\,
            I => \N__1722\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1722\,
            I => \N__1717\
        );

    \I__238\ : InMux
    port map (
            O => \N__1721\,
            I => \N__1712\
        );

    \I__237\ : InMux
    port map (
            O => \N__1720\,
            I => \N__1712\
        );

    \I__236\ : Odrv4
    port map (
            O => \N__1717\,
            I => \arse.seqcounterZ0Z_4\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1712\,
            I => \arse.seqcounterZ0Z_4\
        );

    \I__234\ : CascadeMux
    port map (
            O => \N__1707\,
            I => \N__1703\
        );

    \I__233\ : InMux
    port map (
            O => \N__1706\,
            I => \N__1700\
        );

    \I__232\ : InMux
    port map (
            O => \N__1703\,
            I => \N__1697\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1700\,
            I => \arse.seqcounter_i_4\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__1697\,
            I => \arse.seqcounter_i_4\
        );

    \I__229\ : InMux
    port map (
            O => \N__1692\,
            I => \arses.un2_counter_cry_1\
        );

    \I__228\ : InMux
    port map (
            O => \N__1689\,
            I => \arses.un2_counter_cry_2\
        );

    \I__227\ : InMux
    port map (
            O => \N__1686\,
            I => \arses.un2_counter_cry_3\
        );

    \I__226\ : InMux
    port map (
            O => \N__1683\,
            I => \N__1679\
        );

    \I__225\ : InMux
    port map (
            O => \N__1682\,
            I => \N__1676\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1679\,
            I => \arses.counterZ0Z_5\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1676\,
            I => \arses.counterZ0Z_5\
        );

    \I__222\ : InMux
    port map (
            O => \N__1671\,
            I => \arses.un2_counter_cry_4\
        );

    \I__221\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1664\
        );

    \I__220\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1661\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1664\,
            I => \arses.counterZ0Z_6\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1661\,
            I => \arses.counterZ0Z_6\
        );

    \I__217\ : InMux
    port map (
            O => \N__1656\,
            I => \arses.un2_counter_cry_5\
        );

    \I__216\ : InMux
    port map (
            O => \N__1653\,
            I => \N__1649\
        );

    \I__215\ : InMux
    port map (
            O => \N__1652\,
            I => \N__1646\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1649\,
            I => \arses.counterZ0Z_7\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1646\,
            I => \arses.counterZ0Z_7\
        );

    \I__212\ : InMux
    port map (
            O => \N__1641\,
            I => \arses.un2_counter_cry_6\
        );

    \I__211\ : CascadeMux
    port map (
            O => \N__1638\,
            I => \arse.divseven.N_65_i_cascade_\
        );

    \I__210\ : CascadeMux
    port map (
            O => \N__1635\,
            I => \N__1626\
        );

    \I__209\ : InMux
    port map (
            O => \N__1634\,
            I => \N__1623\
        );

    \I__208\ : InMux
    port map (
            O => \N__1633\,
            I => \N__1620\
        );

    \I__207\ : InMux
    port map (
            O => \N__1632\,
            I => \N__1617\
        );

    \I__206\ : InMux
    port map (
            O => \N__1631\,
            I => \N__1614\
        );

    \I__205\ : InMux
    port map (
            O => \N__1630\,
            I => \N__1607\
        );

    \I__204\ : InMux
    port map (
            O => \N__1629\,
            I => \N__1607\
        );

    \I__203\ : InMux
    port map (
            O => \N__1626\,
            I => \N__1607\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1623\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1620\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1617\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1614\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1607\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__197\ : IoInMux
    port map (
            O => \N__1596\,
            I => \N__1593\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1593\,
            I => \N__1590\
        );

    \I__195\ : Odrv12
    port map (
            O => \N__1590\,
            I => \arse.divseven.doutZ0Z_0\
        );

    \I__194\ : CEMux
    port map (
            O => \N__1587\,
            I => \N__1583\
        );

    \I__193\ : CEMux
    port map (
            O => \N__1586\,
            I => \N__1580\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__1583\,
            I => \N__1577\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1580\,
            I => \N__1574\
        );

    \I__190\ : Span4Mux_h
    port map (
            O => \N__1577\,
            I => \N__1569\
        );

    \I__189\ : Span4Mux_s3_v
    port map (
            O => \N__1574\,
            I => \N__1569\
        );

    \I__188\ : Odrv4
    port map (
            O => \N__1569\,
            I => \arse.divseven.N_65_i_0\
        );

    \I__187\ : InMux
    port map (
            O => \N__1566\,
            I => \N__1563\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1563\,
            I => \arse.seqcounterZ0Z_0\
        );

    \I__185\ : InMux
    port map (
            O => \N__1560\,
            I => \N__1557\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1557\,
            I => \arse.seqcounterZ0Z_1\
        );

    \I__183\ : InMux
    port map (
            O => \N__1554\,
            I => \arse.un1_seqcounter_1_cry_0\
        );

    \I__182\ : InMux
    port map (
            O => \N__1551\,
            I => \N__1548\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1548\,
            I => \arse.seqcounterZ0Z_2\
        );

    \I__180\ : InMux
    port map (
            O => \N__1545\,
            I => \arse.un1_seqcounter_1_cry_1\
        );

    \I__179\ : InMux
    port map (
            O => \N__1542\,
            I => \N__1539\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1539\,
            I => \arse.seqcounterZ1Z_3\
        );

    \I__177\ : InMux
    port map (
            O => \N__1536\,
            I => \arse.un1_seqcounter_1_cry_2\
        );

    \I__176\ : InMux
    port map (
            O => \N__1533\,
            I => \arse.un1_seqcounter_1_cry_3\
        );

    \I__175\ : CascadeMux
    port map (
            O => \N__1530\,
            I => \arse.divseven.N_60_i_cascade_\
        );

    \I__174\ : CEMux
    port map (
            O => \N__1527\,
            I => \N__1524\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1524\,
            I => \N__1521\
        );

    \I__172\ : Odrv12
    port map (
            O => \N__1521\,
            I => \arse.divseven.counter_6_sqmuxa\
        );

    \I__171\ : CascadeMux
    port map (
            O => \N__1518\,
            I => \arse.divseven.N_6_cascade_\
        );

    \I__170\ : CascadeMux
    port map (
            O => \N__1515\,
            I => \arse.divseven.un1_dout_2_sqmuxa_i_o2_0_cascade_\
        );

    \I__169\ : CascadeMux
    port map (
            O => \N__1512\,
            I => \arse.divseven.N_10_cascade_\
        );

    \I__168\ : InMux
    port map (
            O => \N__1509\,
            I => \N__1504\
        );

    \I__167\ : InMux
    port map (
            O => \N__1508\,
            I => \N__1501\
        );

    \I__166\ : InMux
    port map (
            O => \N__1507\,
            I => \N__1495\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1504\,
            I => \N__1490\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1501\,
            I => \N__1490\
        );

    \I__163\ : InMux
    port map (
            O => \N__1500\,
            I => \N__1487\
        );

    \I__162\ : InMux
    port map (
            O => \N__1499\,
            I => \N__1482\
        );

    \I__161\ : InMux
    port map (
            O => \N__1498\,
            I => \N__1482\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1495\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__159\ : Odrv4
    port map (
            O => \N__1490\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1487\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1482\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__156\ : InMux
    port map (
            O => \N__1473\,
            I => \N__1465\
        );

    \I__155\ : InMux
    port map (
            O => \N__1472\,
            I => \N__1462\
        );

    \I__154\ : InMux
    port map (
            O => \N__1471\,
            I => \N__1459\
        );

    \I__153\ : InMux
    port map (
            O => \N__1470\,
            I => \N__1452\
        );

    \I__152\ : InMux
    port map (
            O => \N__1469\,
            I => \N__1452\
        );

    \I__151\ : InMux
    port map (
            O => \N__1468\,
            I => \N__1452\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1465\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__1462\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1459\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1452\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__146\ : CascadeMux
    port map (
            O => \N__1443\,
            I => \N__1439\
        );

    \I__145\ : CascadeMux
    port map (
            O => \N__1442\,
            I => \N__1436\
        );

    \I__144\ : InMux
    port map (
            O => \N__1439\,
            I => \N__1432\
        );

    \I__143\ : InMux
    port map (
            O => \N__1436\,
            I => \N__1429\
        );

    \I__142\ : CascadeMux
    port map (
            O => \N__1435\,
            I => \N__1426\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1432\,
            I => \N__1418\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1429\,
            I => \N__1418\
        );

    \I__139\ : InMux
    port map (
            O => \N__1426\,
            I => \N__1415\
        );

    \I__138\ : InMux
    port map (
            O => \N__1425\,
            I => \N__1412\
        );

    \I__137\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1407\
        );

    \I__136\ : InMux
    port map (
            O => \N__1423\,
            I => \N__1407\
        );

    \I__135\ : Odrv4
    port map (
            O => \N__1418\,
            I => \arse.divseven.sevenZ0\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__1415\,
            I => \arse.divseven.sevenZ0\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1412\,
            I => \arse.divseven.sevenZ0\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__1407\,
            I => \arse.divseven.sevenZ0\
        );

    \I__131\ : IoInMux
    port map (
            O => \N__1398\,
            I => \N__1395\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__1395\,
            I => \N__1392\
        );

    \I__129\ : Odrv12
    port map (
            O => \N__1392\,
            I => \arse.divseven.doutZ0Z_1\
        );

    \I__128\ : IoInMux
    port map (
            O => \N__1389\,
            I => \N__1386\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1386\,
            I => \N__1383\
        );

    \I__126\ : IoSpan4Mux
    port map (
            O => \N__1383\,
            I => \N__1380\
        );

    \I__125\ : Span4Mux_s3_h
    port map (
            O => \N__1380\,
            I => \N__1377\
        );

    \I__124\ : Sp12to4
    port map (
            O => \N__1377\,
            I => \N__1374\
        );

    \I__123\ : Span12Mux_v
    port map (
            O => \N__1374\,
            I => \N__1371\
        );

    \I__122\ : Span12Mux_h
    port map (
            O => \N__1371\,
            I => \N__1368\
        );

    \I__121\ : Odrv12
    port map (
            O => \N__1368\,
            I => \top_pll_nrtthrth.PLLOUTCORE_0\
        );

    \INVarse.diveight.dout_0C\ : INV
    port map (
            O => \INVarse.diveight.dout_0C_net\,
            I => \N__2942\
        );

    \INVarse.divseven.dout_nesr_0C\ : INV
    port map (
            O => \INVarse.divseven.dout_nesr_0C_net\,
            I => \N__2940\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \arses.un2_counter_cry_8\,
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_16_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_6_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1389\,
            GLOBALBUFFEROUTPUT => \PLLOUTCORE_0_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \arse.divseven.dout_esr_1_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1634\,
            in1 => \N__1508\,
            in2 => \N__1443\,
            in3 => \N__1473\,
            lcout => \arse.divseven.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2936\,
            ce => \N__1587\,
            sr => \N__2879\
        );

    \arse.divseven.seven_RNO_0_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1425\,
            in2 => \_gnd_net_\,
            in3 => \N__1471\,
            lcout => OPEN,
            ltout => \arse.divseven.N_60_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.seven_RNO_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1632\,
            in1 => \N__1500\,
            in2 => \N__1530\,
            in3 => \N__3130\,
            lcout => \arse.divseven.counter_6_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.seven_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3372\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \arse.divseven.sevenZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2935\,
            ce => \N__1527\,
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_ns_2_0__m5_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110010110011"
        )
    port map (
            in0 => \N__1633\,
            in1 => \N__1509\,
            in2 => \N__1442\,
            in3 => \N__1472\,
            lcout => OPEN,
            ltout => \arse.divseven.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_1_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__3125\,
            in1 => \_gnd_net_\,
            in2 => \N__1518\,
            in3 => \_gnd_net_\,
            lcout => \arse.divseven.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_ns_2_0__m3_s_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__1499\,
            in1 => \N__1424\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \arse.divseven.un1_dout_2_sqmuxa_i_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_0_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010100000000"
        )
    port map (
            in0 => \N__1470\,
            in1 => \N__1630\,
            in2 => \N__1515\,
            in3 => \N__3097\,
            lcout => \arse.divseven.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_ns_2_0__m9_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100111010101"
        )
    port map (
            in0 => \N__1629\,
            in1 => \N__1507\,
            in2 => \N__1435\,
            in3 => \N__1469\,
            lcout => OPEN,
            ltout => \arse.divseven.N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_2_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1512\,
            in3 => \N__3096\,
            lcout => \arse.divseven.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_RNI8ECT_0_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__1498\,
            in1 => \N__1468\,
            in2 => \N__1635\,
            in3 => \N__1423\,
            lcout => OPEN,
            ltout => \arse.divseven.N_65_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_RNI04101_0_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1638\,
            in3 => \N__2841\,
            lcout => \arse.divseven.N_65_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_nesr_0_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1631\,
            lcout => \arse.divseven.doutZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.divseven.dout_nesr_0C_net\,
            ce => \N__1586\,
            sr => \N__2842\
        );

    \arse.seqreset_e_0_RNIOLK2_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3074\,
            lcout => \arse.seqreset_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqreset_e_0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1725\,
            lcout => \arse.seqresetZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2938\,
            ce => \N__2325\,
            sr => \_gnd_net_\
        );

    \arse.seqcounter_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2307\,
            in1 => \N__1566\,
            in2 => \N__1707\,
            in3 => \N__1706\,
            lcout => \arse.seqcounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \arse.un1_seqcounter_1_cry_0\,
            clk => \N__2934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqcounter_1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2309\,
            in1 => \N__1560\,
            in2 => \_gnd_net_\,
            in3 => \N__1554\,
            lcout => \arse.seqcounterZ0Z_1\,
            ltout => OPEN,
            carryin => \arse.un1_seqcounter_1_cry_0\,
            carryout => \arse.un1_seqcounter_1_cry_1\,
            clk => \N__2934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqcounter_2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2308\,
            in1 => \N__1551\,
            in2 => \_gnd_net_\,
            in3 => \N__1545\,
            lcout => \arse.seqcounterZ0Z_2\,
            ltout => OPEN,
            carryin => \arse.un1_seqcounter_1_cry_1\,
            carryout => \arse.un1_seqcounter_1_cry_2\,
            clk => \N__2934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqcounter_3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2310\,
            in1 => \N__1542\,
            in2 => \_gnd_net_\,
            in3 => \N__1536\,
            lcout => \arse.seqcounterZ1Z_3\,
            ltout => OPEN,
            carryin => \arse.un1_seqcounter_1_cry_2\,
            carryout => \arse.un1_seqcounter_1_cry_3\,
            clk => \N__2934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqcounter_4_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__1721\,
            in1 => \N__2311\,
            in2 => \_gnd_net_\,
            in3 => \N__1533\,
            lcout => \arse.seqcounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2934\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqcounter_RNIEP0A_4_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1720\,
            lcout => \arse.seqcounter_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIA58_5_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1652\,
            in1 => \N__1667\,
            in2 => \N__1782\,
            in3 => \N__1682\,
            lcout => \arses.un1_counterlto8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.un2_counter_cry_1_c_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1896\,
            in2 => \N__1875\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \arses.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_2_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2201\,
            in1 => \N__1932\,
            in2 => \_gnd_net_\,
            in3 => \N__1692\,
            lcout => \arses.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_1\,
            carryout => \arses.un2_counter_cry_2\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_3_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2193\,
            in1 => \N__1944\,
            in2 => \_gnd_net_\,
            in3 => \N__1689\,
            lcout => \arses.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_2\,
            carryout => \arses.un2_counter_cry_3\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_4_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2202\,
            in1 => \N__1919\,
            in2 => \_gnd_net_\,
            in3 => \N__1686\,
            lcout => \arses.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_3\,
            carryout => \arses.un2_counter_cry_4\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_5_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2194\,
            in1 => \N__1683\,
            in2 => \_gnd_net_\,
            in3 => \N__1671\,
            lcout => \arses.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_4\,
            carryout => \arses.un2_counter_cry_5\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_6_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2203\,
            in1 => \N__1668\,
            in2 => \_gnd_net_\,
            in3 => \N__1656\,
            lcout => \arses.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_5\,
            carryout => \arses.un2_counter_cry_6\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_7_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2195\,
            in1 => \N__1653\,
            in2 => \_gnd_net_\,
            in3 => \N__1641\,
            lcout => \arses.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_6\,
            carryout => \arses.un2_counter_cry_7\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_8_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2204\,
            in1 => \N__1781\,
            in2 => \_gnd_net_\,
            in3 => \N__1767\,
            lcout => \arses.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_7\,
            carryout => \arses.un2_counter_cry_8\,
            clk => \N__2473\,
            ce => 'H',
            sr => \N__1852\
        );

    \arses.counter_9_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2192\,
            in1 => \N__1794\,
            in2 => \_gnd_net_\,
            in3 => \N__1764\,
            lcout => \arses.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \arses.un2_counter_cry_9\,
            clk => \N__2474\,
            ce => 'H',
            sr => \N__1854\
        );

    \arses.counter_10_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2198\,
            in1 => \N__1827\,
            in2 => \_gnd_net_\,
            in3 => \N__1761\,
            lcout => \arses.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_9\,
            carryout => \arses.un2_counter_cry_10\,
            clk => \N__2474\,
            ce => 'H',
            sr => \N__1854\
        );

    \arses.counter_11_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2190\,
            in1 => \N__1808\,
            in2 => \_gnd_net_\,
            in3 => \N__1758\,
            lcout => \arses.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_10\,
            carryout => \arses.un2_counter_cry_11\,
            clk => \N__2474\,
            ce => 'H',
            sr => \N__1854\
        );

    \arses.counter_12_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2199\,
            in1 => \N__2040\,
            in2 => \_gnd_net_\,
            in3 => \N__1755\,
            lcout => \arses.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_11\,
            carryout => \arses.un2_counter_cry_12\,
            clk => \N__2474\,
            ce => 'H',
            sr => \N__1854\
        );

    \arses.counter_13_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2191\,
            in1 => \N__2055\,
            in2 => \_gnd_net_\,
            in3 => \N__1752\,
            lcout => \arses.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_12\,
            carryout => \arses.un2_counter_cry_13\,
            clk => \N__2474\,
            ce => 'H',
            sr => \N__1854\
        );

    \arses.counter_14_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2200\,
            in1 => \N__2067\,
            in2 => \_gnd_net_\,
            in3 => \N__1749\,
            lcout => \arses.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2474\,
            ce => 'H',
            sr => \N__1854\
        );

    \masterreset_ibuf_RNIKP26_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => masterreset_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_0_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2981\,
            lcout => \arse.diveight.doutZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.diveight.dout_0C_net\,
            ce => 'H',
            sr => \N__2887\
        );

    \arse.diveight.counter_2_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110000000000"
        )
    port map (
            in0 => \N__1961\,
            in1 => \N__2977\,
            in2 => \N__1974\,
            in3 => \N__3139\,
            lcout => \arse.diveight.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_1_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3137\,
            in2 => \N__1962\,
            in3 => \N__1970\,
            lcout => \arse.diveight.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_0_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__3138\,
            in1 => \N__1957\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \arse.diveight.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI1L5_2_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__1943\,
            in1 => \N__1931\,
            in2 => \_gnd_net_\,
            in3 => \N__1890\,
            lcout => OPEN,
            ltout => \arses.un1_counterlto4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOKH_1_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__1920\,
            in1 => \N__1867\,
            in2 => \N__1905\,
            in3 => \N__1902\,
            lcout => \arses.un1_counterlt11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_0_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__1891\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2197\,
            lcout => \arses.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2471\,
            ce => 'H',
            sr => \N__1853\
        );

    \arses.counter_1_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__2196\,
            in1 => \_gnd_net_\,
            in2 => \N__1874\,
            in3 => \N__1892\,
            lcout => \arses.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2471\,
            ce => 'H',
            sr => \N__1853\
        );

    \arses.counter_RNI04C4_9_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1826\,
            in1 => \N__1815\,
            in2 => \N__1809\,
            in3 => \N__1793\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOS0A_14_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__2066\,
            in1 => \N__2054\,
            in2 => \N__2043\,
            in3 => \N__2039\,
            lcout => \arses.counter8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_4_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__2552\,
            in1 => \N__2358\,
            in2 => \N__2598\,
            in3 => \N__2375\,
            lcout => \debounceconsolereset.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_2_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__2550\,
            in1 => \N__2007\,
            in2 => \N__2028\,
            in3 => \N__2596\,
            lcout => \debounceconsolereset.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_RNO_1_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2024\,
            in1 => \N__2374\,
            in2 => \N__1997\,
            in3 => \N__2520\,
            lcout => \debounceconsolereset.out_cnv_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNISLFD_2_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2373\,
            in1 => \N__1989\,
            in2 => \_gnd_net_\,
            in3 => \N__2023\,
            lcout => \debounceconsolereset.un1_counterlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_3_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__2551\,
            in1 => \N__2385\,
            in2 => \N__1998\,
            in3 => \N__2597\,
            lcout => \debounceconsolereset.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_0_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__2521\,
            in1 => \N__2591\,
            in2 => \_gnd_net_\,
            in3 => \N__2553\,
            lcout => \debounceconsolereset.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_1_c_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2491\,
            in2 => \N__2525\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \debounceconsolereset.un3_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2022\,
            in2 => \_gnd_net_\,
            in3 => \N__2001\,
            lcout => \debounceconsolereset.un3_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_1\,
            carryout => \debounceconsolereset.un3_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1996\,
            in2 => \_gnd_net_\,
            in3 => \N__2379\,
            lcout => \debounceconsolereset.un3_counter_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_2\,
            carryout => \debounceconsolereset.un3_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_3_THRU_LUT4_0_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2376\,
            in2 => \_gnd_net_\,
            in3 => \N__2352\,
            lcout => \debounceconsolereset.un3_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_3\,
            carryout => \debounceconsolereset.un3_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_4_THRU_LUT4_0_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2110\,
            in2 => \_gnd_net_\,
            in3 => \N__2349\,
            lcout => \debounceconsolereset.un3_counter_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_4\,
            carryout => \debounceconsolereset.un3_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_6_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__2085\,
            in1 => \N__2595\,
            in2 => \N__2559\,
            in3 => \N__2346\,
            lcout => \debounceconsolereset.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__2334\,
            in1 => \N__2132\,
            in2 => \_gnd_net_\,
            in3 => \N__2189\,
            lcout => \clock_out_RNIR6ER\,
            ltout => \clock_out_RNIR6ER_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNI4RTH1_6_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__2109\,
            in1 => \N__2083\,
            in2 => \N__2343\,
            in3 => \N__2340\,
            lcout => \debounceconsolereset.counter_RNI4RTH1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2333\,
            in1 => \N__2133\,
            in2 => \_gnd_net_\,
            in3 => \N__2205\,
            lcout => \arses.clock_out_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_5_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__2554\,
            in1 => \N__2112\,
            in2 => \N__2121\,
            in3 => \N__2590\,
            lcout => \debounceconsolereset.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_RNO_0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__2111\,
            in1 => \N__2094\,
            in2 => \N__2498\,
            in3 => \N__2084\,
            lcout => OPEN,
            ltout => \debounceconsolereset.out_cnv_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__2616\,
            in1 => \N__2589\,
            in2 => \N__2601\,
            in3 => \N__3239\,
            lcout => apureset_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_1_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__2588\,
            in1 => \N__2555\,
            in2 => \N__2499\,
            in3 => \N__2526\,
            lcout => \debounceconsolereset.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2472\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.counter_1_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__2726\,
            in1 => \N__2433\,
            in2 => \N__2409\,
            in3 => \N__2670\,
            lcout => \arse.arse.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2943\,
            ce => 'H',
            sr => \N__2866\
        );

    \arse.arse.counter_2_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__2727\,
            in1 => \N__2810\,
            in2 => \N__2787\,
            in3 => \N__2671\,
            lcout => \arse.arse.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2943\,
            ce => 'H',
            sr => \N__2866\
        );

    \arse.arse.counter_RNIHKTF1_1_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__2808\,
            in1 => \N__2401\,
            in2 => \_gnd_net_\,
            in3 => \N__2430\,
            lcout => \arse.un1_counterlt4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2478\,
            lcout => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.counter_0_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__2811\,
            in1 => \N__2716\,
            in2 => \_gnd_net_\,
            in3 => \N__2432\,
            lcout => \arse.arse.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2945\,
            ce => 'H',
            sr => \N__2880\
        );

    \arse.arse.counter_3_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__2717\,
            in1 => \N__2748\,
            in2 => \N__2775\,
            in3 => \N__2675\,
            lcout => \arse.arse.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2945\,
            ce => 'H',
            sr => \N__2880\
        );

    \arse.arse.un16_counter_cry_1_c_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2431\,
            in2 => \N__2408\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_6_0_\,
            carryout => \arse.arse.un16_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.un16_counter_cry_1_THRU_LUT4_0_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2809\,
            in2 => \_gnd_net_\,
            in3 => \N__2778\,
            lcout => \arse.arse.un16_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \arse.arse.un16_counter_cry_1\,
            carryout => \arse.arse.un16_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.un16_counter_cry_2_THRU_LUT4_0_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2747\,
            in2 => \_gnd_net_\,
            in3 => \N__2766\,
            lcout => \arse.arse.un16_counter_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \arse.arse.un16_counter_cry_2\,
            carryout => \arse.arse.un16_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.counter_4_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__2760\,
            in1 => \N__2715\,
            in2 => \N__2682\,
            in3 => \N__2763\,
            lcout => \arse.arse.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2944\,
            ce => 'H',
            sr => \N__2888\
        );

    \arse.arse.counter_RNIRIUV_4_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2759\,
            in2 => \_gnd_net_\,
            in3 => \N__2746\,
            lcout => \arse.un1_counterlto4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.ddd.Q_esr_RNO_LC_18_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3284\,
            in2 => \_gnd_net_\,
            in3 => \N__2622\,
            lcout => \arse.ddd.N_33_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.clock_out_RNIM09F_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3269\,
            in2 => \_gnd_net_\,
            in3 => \N__2632\,
            lcout => OPEN,
            ltout => \arse.G_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.seqreset_e_0_RNIQTP13_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2713\,
            in1 => \N__2677\,
            in2 => \N__2730\,
            in3 => \N__3127\,
            lcout => \arse.seqreset_e_0_RNIQTPZ0Z13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.arse.clock_out_LC_18_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__2714\,
            in1 => \N__2678\,
            in2 => \N__2640\,
            in3 => \N__3128\,
            lcout => \arse.clock_out_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2946\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.ddd.Q_esr_RNO_0_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__2712\,
            in1 => \N__2676\,
            in2 => \N__2639\,
            in3 => \N__3126\,
            lcout => \arse.ddd.Q_esr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.ddd.Q_esr_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__3255\,
            in1 => \N__3218\,
            in2 => \N__3146\,
            in3 => \N__3206\,
            lcout => cpureset_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2947\,
            ce => \N__3297\,
            sr => \N__3291\
        );

    \arse.l2.un1_Q_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__3219\,
            in1 => \N__3207\,
            in2 => \N__3273\,
            in3 => \N__3129\,
            lcout => \G_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.l1.N_23_0_i_LC_20_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__3036\,
            in1 => \N__3199\,
            in2 => \N__3164\,
            in3 => \N__3147\,
            lcout => \G_74\,
            ltout => \G_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.io_0_RNIIG08_LC_20_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__3030\,
            in1 => \_gnd_net_\,
            in2 => \N__3018\,
            in3 => \_gnd_net_\,
            lcout => arse_un1_apuclk_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_1_LC_30_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2994\,
            lcout => \arse.diveight.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2948\,
            ce => 'H',
            sr => \N__2892\
        );
end \INTERFACE\;
