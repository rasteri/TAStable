// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 8 2024 23:35:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    led5,
    lcol2,
    led6,
    led2,
    lcol1,
    cpuclk,
    apureset,
    led7,
    led3,
    lcol4,
    cpureset,
    apusync,
    PACKAGEPIN,
    masterreset,
    led8,
    led4,
    lcol3,
    led1,
    consolereset,
    apuclk);

    output led5;
    output lcol2;
    output led6;
    output led2;
    output lcol1;
    output cpuclk;
    output apureset;
    output led7;
    output led3;
    output lcol4;
    output cpureset;
    input apusync;
    input PACKAGEPIN;
    input masterreset;
    output led8;
    output led4;
    output lcol3;
    output led1;
    input consolereset;
    output apuclk;

    wire N__3600;
    wire N__3599;
    wire N__3598;
    wire N__3589;
    wire N__3588;
    wire N__3587;
    wire N__3580;
    wire N__3579;
    wire N__3578;
    wire N__3571;
    wire N__3570;
    wire N__3569;
    wire N__3562;
    wire N__3561;
    wire N__3560;
    wire N__3553;
    wire N__3552;
    wire N__3551;
    wire N__3544;
    wire N__3543;
    wire N__3542;
    wire N__3535;
    wire N__3534;
    wire N__3533;
    wire N__3526;
    wire N__3525;
    wire N__3524;
    wire N__3517;
    wire N__3516;
    wire N__3515;
    wire N__3508;
    wire N__3507;
    wire N__3506;
    wire N__3499;
    wire N__3498;
    wire N__3497;
    wire N__3490;
    wire N__3489;
    wire N__3488;
    wire N__3481;
    wire N__3480;
    wire N__3479;
    wire N__3472;
    wire N__3471;
    wire N__3470;
    wire N__3463;
    wire N__3462;
    wire N__3461;
    wire N__3454;
    wire N__3453;
    wire N__3452;
    wire N__3445;
    wire N__3444;
    wire N__3443;
    wire N__3436;
    wire N__3435;
    wire N__3434;
    wire N__3427;
    wire N__3426;
    wire N__3425;
    wire N__3418;
    wire N__3417;
    wire N__3416;
    wire N__3399;
    wire N__3398;
    wire N__3395;
    wire N__3394;
    wire N__3391;
    wire N__3390;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3372;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3344;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3330;
    wire N__3327;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3302;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3273;
    wire N__3270;
    wire N__3269;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3239;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3219;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3207;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3199;
    wire N__3194;
    wire N__3191;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3147;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3139;
    wire N__3138;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3130;
    wire N__3129;
    wire N__3128;
    wire N__3127;
    wire N__3126;
    wire N__3125;
    wire N__3122;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3098;
    wire N__3097;
    wire N__3096;
    wire N__3093;
    wire N__3088;
    wire N__3083;
    wire N__3080;
    wire N__3075;
    wire N__3074;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2981;
    wire N__2978;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2948;
    wire N__2947;
    wire N__2946;
    wire N__2945;
    wire N__2944;
    wire N__2943;
    wire N__2942;
    wire N__2941;
    wire N__2940;
    wire N__2939;
    wire N__2938;
    wire N__2937;
    wire N__2936;
    wire N__2935;
    wire N__2934;
    wire N__2933;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2888;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2880;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2842;
    wire N__2841;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2811;
    wire N__2810;
    wire N__2809;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2748;
    wire N__2747;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2730;
    wire N__2727;
    wire N__2726;
    wire N__2721;
    wire N__2718;
    wire N__2717;
    wire N__2716;
    wire N__2715;
    wire N__2714;
    wire N__2713;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2693;
    wire N__2682;
    wire N__2679;
    wire N__2678;
    wire N__2677;
    wire N__2676;
    wire N__2675;
    wire N__2672;
    wire N__2671;
    wire N__2670;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2652;
    wire N__2649;
    wire N__2640;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2632;
    wire N__2625;
    wire N__2622;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2597;
    wire N__2596;
    wire N__2595;
    wire N__2592;
    wire N__2591;
    wire N__2590;
    wire N__2589;
    wire N__2588;
    wire N__2583;
    wire N__2580;
    wire N__2575;
    wire N__2568;
    wire N__2559;
    wire N__2556;
    wire N__2555;
    wire N__2554;
    wire N__2553;
    wire N__2552;
    wire N__2551;
    wire N__2550;
    wire N__2547;
    wire N__2542;
    wire N__2533;
    wire N__2526;
    wire N__2525;
    wire N__2522;
    wire N__2521;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2509;
    wire N__2506;
    wire N__2499;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2491;
    wire N__2486;
    wire N__2483;
    wire N__2478;
    wire N__2475;
    wire N__2474;
    wire N__2473;
    wire N__2472;
    wire N__2471;
    wire N__2470;
    wire N__2469;
    wire N__2466;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2432;
    wire N__2431;
    wire N__2430;
    wire N__2427;
    wire N__2424;
    wire N__2421;
    wire N__2418;
    wire N__2409;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2401;
    wire N__2398;
    wire N__2395;
    wire N__2392;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2376;
    wire N__2375;
    wire N__2374;
    wire N__2373;
    wire N__2370;
    wire N__2363;
    wire N__2358;
    wire N__2355;
    wire N__2352;
    wire N__2349;
    wire N__2346;
    wire N__2343;
    wire N__2340;
    wire N__2337;
    wire N__2334;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2326;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2311;
    wire N__2310;
    wire N__2309;
    wire N__2308;
    wire N__2307;
    wire N__2304;
    wire N__2301;
    wire N__2298;
    wire N__2295;
    wire N__2292;
    wire N__2285;
    wire N__2280;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2262;
    wire N__2257;
    wire N__2254;
    wire N__2251;
    wire N__2248;
    wire N__2245;
    wire N__2242;
    wire N__2239;
    wire N__2236;
    wire N__2233;
    wire N__2230;
    wire N__2227;
    wire N__2224;
    wire N__2221;
    wire N__2218;
    wire N__2215;
    wire N__2212;
    wire N__2205;
    wire N__2204;
    wire N__2203;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2196;
    wire N__2195;
    wire N__2194;
    wire N__2193;
    wire N__2192;
    wire N__2191;
    wire N__2190;
    wire N__2189;
    wire N__2186;
    wire N__2177;
    wire N__2170;
    wire N__2165;
    wire N__2158;
    wire N__2151;
    wire N__2148;
    wire N__2133;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2121;
    wire N__2118;
    wire N__2115;
    wire N__2112;
    wire N__2111;
    wire N__2110;
    wire N__2109;
    wire N__2104;
    wire N__2099;
    wire N__2094;
    wire N__2091;
    wire N__2088;
    wire N__2085;
    wire N__2084;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2067;
    wire N__2066;
    wire N__2063;
    wire N__2060;
    wire N__2055;
    wire N__2054;
    wire N__2051;
    wire N__2048;
    wire N__2043;
    wire N__2040;
    wire N__2039;
    wire N__2036;
    wire N__2033;
    wire N__2028;
    wire N__2025;
    wire N__2024;
    wire N__2023;
    wire N__2022;
    wire N__2015;
    wire N__2012;
    wire N__2007;
    wire N__2004;
    wire N__2001;
    wire N__1998;
    wire N__1997;
    wire N__1996;
    wire N__1993;
    wire N__1990;
    wire N__1989;
    wire N__1986;
    wire N__1979;
    wire N__1974;
    wire N__1971;
    wire N__1970;
    wire N__1965;
    wire N__1962;
    wire N__1961;
    wire N__1958;
    wire N__1957;
    wire N__1954;
    wire N__1949;
    wire N__1944;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1932;
    wire N__1931;
    wire N__1928;
    wire N__1925;
    wire N__1920;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1905;
    wire N__1902;
    wire N__1899;
    wire N__1896;
    wire N__1893;
    wire N__1892;
    wire N__1891;
    wire N__1890;
    wire N__1887;
    wire N__1880;
    wire N__1875;
    wire N__1874;
    wire N__1871;
    wire N__1868;
    wire N__1867;
    wire N__1864;
    wire N__1859;
    wire N__1854;
    wire N__1853;
    wire N__1852;
    wire N__1849;
    wire N__1846;
    wire N__1843;
    wire N__1840;
    wire N__1835;
    wire N__1832;
    wire N__1827;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1815;
    wire N__1812;
    wire N__1809;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1794;
    wire N__1793;
    wire N__1790;
    wire N__1787;
    wire N__1782;
    wire N__1781;
    wire N__1778;
    wire N__1775;
    wire N__1772;
    wire N__1767;
    wire N__1764;
    wire N__1761;
    wire N__1758;
    wire N__1755;
    wire N__1752;
    wire N__1749;
    wire N__1746;
    wire N__1743;
    wire N__1740;
    wire N__1737;
    wire N__1734;
    wire N__1731;
    wire N__1728;
    wire N__1725;
    wire N__1722;
    wire N__1721;
    wire N__1720;
    wire N__1717;
    wire N__1712;
    wire N__1707;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1697;
    wire N__1692;
    wire N__1689;
    wire N__1686;
    wire N__1683;
    wire N__1682;
    wire N__1679;
    wire N__1676;
    wire N__1671;
    wire N__1668;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1656;
    wire N__1653;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1641;
    wire N__1638;
    wire N__1635;
    wire N__1634;
    wire N__1633;
    wire N__1632;
    wire N__1631;
    wire N__1630;
    wire N__1629;
    wire N__1626;
    wire N__1623;
    wire N__1620;
    wire N__1617;
    wire N__1614;
    wire N__1607;
    wire N__1596;
    wire N__1593;
    wire N__1590;
    wire N__1587;
    wire N__1586;
    wire N__1583;
    wire N__1580;
    wire N__1577;
    wire N__1574;
    wire N__1569;
    wire N__1566;
    wire N__1563;
    wire N__1560;
    wire N__1557;
    wire N__1554;
    wire N__1551;
    wire N__1548;
    wire N__1545;
    wire N__1542;
    wire N__1539;
    wire N__1536;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1524;
    wire N__1521;
    wire N__1518;
    wire N__1515;
    wire N__1512;
    wire N__1509;
    wire N__1508;
    wire N__1507;
    wire N__1504;
    wire N__1501;
    wire N__1500;
    wire N__1499;
    wire N__1498;
    wire N__1495;
    wire N__1490;
    wire N__1487;
    wire N__1482;
    wire N__1473;
    wire N__1472;
    wire N__1471;
    wire N__1470;
    wire N__1469;
    wire N__1468;
    wire N__1465;
    wire N__1462;
    wire N__1459;
    wire N__1452;
    wire N__1443;
    wire N__1442;
    wire N__1439;
    wire N__1436;
    wire N__1435;
    wire N__1432;
    wire N__1429;
    wire N__1426;
    wire N__1425;
    wire N__1424;
    wire N__1423;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1407;
    wire N__1398;
    wire N__1395;
    wire N__1392;
    wire N__1389;
    wire N__1386;
    wire N__1383;
    wire N__1380;
    wire N__1377;
    wire N__1374;
    wire N__1371;
    wire N__1368;
    wire \top_pll_nrtthrth.PLLOUTCORE_0 ;
    wire GNDG0;
    wire VCCG0;
    wire \arse.divseven.doutZ0Z_1 ;
    wire \arse.divseven.N_60_i_cascade_ ;
    wire \arse.divseven.counter_6_sqmuxa ;
    wire \arse.divseven.N_6_cascade_ ;
    wire \arse.divseven.un1_dout_2_sqmuxa_i_o2_0_cascade_ ;
    wire \arse.divseven.N_10_cascade_ ;
    wire \arse.divseven.counterZ0Z_1 ;
    wire \arse.divseven.counterZ0Z_0 ;
    wire \arse.divseven.sevenZ0 ;
    wire \arse.divseven.N_65_i_cascade_ ;
    wire \arse.divseven.counterZ0Z_2 ;
    wire \arse.divseven.doutZ0Z_0 ;
    wire \INVarse.divseven.dout_nesr_0C_net ;
    wire \arse.divseven.N_65_i_0 ;
    wire \arse.seqcounterZ0Z_0 ;
    wire bfn_6_9_0_;
    wire \arse.seqcounterZ0Z_1 ;
    wire \arse.un1_seqcounter_1_cry_0 ;
    wire \arse.seqcounterZ0Z_2 ;
    wire \arse.un1_seqcounter_1_cry_1 ;
    wire \arse.seqcounterZ1Z_3 ;
    wire \arse.un1_seqcounter_1_cry_2 ;
    wire \arse.un1_seqcounter_1_cry_3 ;
    wire \arse.seqcounterZ0Z_4 ;
    wire \arse.seqcounter_i_4 ;
    wire bfn_9_4_0_;
    wire \arses.un2_counter_cry_1 ;
    wire \arses.un2_counter_cry_2 ;
    wire \arses.un2_counter_cry_3 ;
    wire \arses.counterZ0Z_5 ;
    wire \arses.un2_counter_cry_4 ;
    wire \arses.counterZ0Z_6 ;
    wire \arses.un2_counter_cry_5 ;
    wire \arses.counterZ0Z_7 ;
    wire \arses.un2_counter_cry_6 ;
    wire \arses.counterZ0Z_8 ;
    wire \arses.un2_counter_cry_7 ;
    wire \arses.un2_counter_cry_8 ;
    wire bfn_9_5_0_;
    wire \arses.un2_counter_cry_9 ;
    wire \arses.un2_counter_cry_10 ;
    wire \arses.un2_counter_cry_11 ;
    wire \arses.un2_counter_cry_12 ;
    wire \arses.un2_counter_cry_13 ;
    wire \arse.diveight.doutZ0Z_0 ;
    wire \INVarse.diveight.dout_0C_net ;
    wire \arse.diveight.counterZ0Z_1 ;
    wire \arse.diveight.counterZ0Z_0 ;
    wire \arses.counterZ0Z_3 ;
    wire \arses.counterZ0Z_2 ;
    wire \arses.counterZ0Z_4 ;
    wire \arses.un1_counterlto4_2_cascade_ ;
    wire \arses.un1_counterlto8_2 ;
    wire \arses.counterZ0Z_0 ;
    wire \arses.counterZ0Z_1 ;
    wire masterreset_c_i;
    wire \arses.counterZ0Z_10 ;
    wire \arses.un1_counterlt11 ;
    wire \arses.counterZ0Z_11 ;
    wire \arses.counterZ0Z_9 ;
    wire \arses.counterZ0Z_14 ;
    wire \arses.counterZ0Z_13 ;
    wire \arses.un1_counterlt13_0_cascade_ ;
    wire \arses.counterZ0Z_12 ;
    wire bfn_11_4_0_;
    wire \debounceconsolereset.counterZ0Z_2 ;
    wire \debounceconsolereset.un3_counter_cry_1_THRU_CO ;
    wire \debounceconsolereset.un3_counter_cry_1 ;
    wire \debounceconsolereset.counterZ0Z_3 ;
    wire \debounceconsolereset.un3_counter_cry_2_THRU_CO ;
    wire \debounceconsolereset.un3_counter_cry_2 ;
    wire \debounceconsolereset.counterZ0Z_4 ;
    wire \debounceconsolereset.un3_counter_cry_3_THRU_CO ;
    wire \debounceconsolereset.un3_counter_cry_3 ;
    wire \debounceconsolereset.un3_counter_cry_4 ;
    wire \debounceconsolereset.un3_counter_cry_5 ;
    wire clock_out_RNIR6ER_cascade_;
    wire \debounceconsolereset.un1_counterlt6 ;
    wire masterreset_c;
    wire \arses.counter8 ;
    wire \arses.clock_out_i ;
    wire \debounceconsolereset.un3_counter_cry_4_THRU_CO ;
    wire \debounceconsolereset.counterZ0Z_5 ;
    wire \debounceconsolereset.out_cnv_3 ;
    wire \debounceconsolereset.counterZ0Z_6 ;
    wire consolereset_c;
    wire \debounceconsolereset.out_cnv_4_cascade_ ;
    wire clock_out_RNIR6ER;
    wire \debounceconsolereset.counter_RNI4RTH1Z0Z_6 ;
    wire \debounceconsolereset.counterZ0Z_0 ;
    wire \debounceconsolereset.counterZ0Z_1 ;
    wire PACKAGEPIN_0_c_g;
    wire GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO;
    wire \arse.arse.counterZ0Z_0 ;
    wire \arse.arse.counterZ0Z_1 ;
    wire bfn_16_6_0_;
    wire \arse.arse.counterZ0Z_2 ;
    wire \arse.arse.un16_counter_cry_1_THRU_CO ;
    wire \arse.arse.un16_counter_cry_1 ;
    wire \arse.arse.un16_counter_cry_2_THRU_CO ;
    wire \arse.arse.un16_counter_cry_2 ;
    wire \arse.arse.un16_counter_cry_3 ;
    wire \arse.arse.counterZ0Z_4 ;
    wire \arse.arse.counterZ0Z_3 ;
    wire \arse.G_2_0_cascade_ ;
    wire \arse.un1_counterlto4_0 ;
    wire \arse.un1_counterlt4 ;
    wire \arse.clock_out_i ;
    wire \arse.ddd.Q_esr_RNOZ0Z_0 ;
    wire CONSTANT_ONE_NET;
    wire \arse.ddd.N_33_0 ;
    wire \arse.seqreset_e_0_RNIQTPZ0Z13 ;
    wire apureset_c;
    wire G_73;
    wire apusync_c;
    wire cpureset_c;
    wire \arse.seqresetZ0 ;
    wire G_74;
    wire \arse.divseven.io_0_D_IN_0 ;
    wire G_74_cascade_;
    wire arse_un1_apuclk_i;
    wire \arse.diveight.counterZ0Z_2 ;
    wire \arse.diveight.doutZ0Z_1 ;
    wire _gnd_net_;
    wire PLLOUTCORE_0_g;
    wire \arse.seqreset_i ;

    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .TEST_MODE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FILTER_RANGE=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_RELATIVE=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVR=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVQ=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVF=7'b0011111;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \top_pll_nrtthrth.top_pll_nrtthrth_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\top_pll_nrtthrth.PLLOUTCORE_0 ),
            .REFERENCECLK(N__2445),
            .RESETB(N__2318),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF PACKAGEPIN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3598),
            .GLOBALBUFFEROUTPUT(PACKAGEPIN_0_c_g));
    IO_PAD PACKAGEPIN_ibuf_gb_io_iopad (
            .OE(N__3600),
            .DIN(N__3599),
            .DOUT(N__3598),
            .PACKAGEPIN(PACKAGEPIN));
    defparam PACKAGEPIN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam PACKAGEPIN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO PACKAGEPIN_ibuf_gb_io_preio (
            .PADOEN(N__3600),
            .PADOUT(N__3599),
            .PADIN(N__3598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol1_obuf_iopad (
            .OE(N__3589),
            .DIN(N__3588),
            .DOUT(N__3587),
            .PACKAGEPIN(lcol1));
    defparam lcol1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol1_obuf_preio (
            .PADOEN(N__3589),
            .PADOUT(N__3588),
            .PADIN(N__3587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD masterreset_ibuf_iopad (
            .OE(N__3580),
            .DIN(N__3579),
            .DOUT(N__3578),
            .PACKAGEPIN(masterreset));
    defparam masterreset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam masterreset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO masterreset_ibuf_preio (
            .PADOEN(N__3580),
            .PADOUT(N__3579),
            .PADIN(N__3578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(masterreset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam cpureset_obuf_iopad.PULLUP=1'b0;
    defparam cpureset_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD cpureset_obuf_iopad (
            .OE(N__3571),
            .DIN(N__3570),
            .DOUT(N__3569),
            .PACKAGEPIN(cpureset));
    defparam cpureset_obuf_preio.NEG_TRIGGER=1'b0;
    defparam cpureset_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO cpureset_obuf_preio (
            .PADOEN(N__3571),
            .PADOUT(N__3570),
            .PADIN(N__3569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3177),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led8_obuft_iopad (
            .OE(N__3562),
            .DIN(N__3561),
            .DOUT(N__3560),
            .PACKAGEPIN(led8));
    defparam led8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led8_obuft_preio (
            .PADOEN(N__3562),
            .PADOUT(N__3561),
            .PADIN(N__3560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.divseven.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.divseven.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.divseven.io_0_iopad  (
            .OE(N__3553),
            .DIN(N__3552),
            .DOUT(N__3551),
            .PACKAGEPIN());
    defparam \arse.divseven.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.divseven.io_0_preio  (
            .PADOEN(N__3553),
            .PADOUT(N__3552),
            .PADIN(N__3551),
            .CLOCKENABLE(),
            .DOUT1(N__1398),
            .OUTPUTENABLE(N__3389),
            .DIN0(\arse.divseven.io_0_D_IN_0 ),
            .DOUT0(N__1596),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__2933));
    IO_PAD lcol3_obuf_iopad (
            .OE(N__3544),
            .DIN(N__3543),
            .DOUT(N__3542),
            .PACKAGEPIN(lcol3));
    defparam lcol3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol3_obuf_preio (
            .PADOEN(N__3544),
            .PADOUT(N__3543),
            .PADIN(N__3542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3379),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam apuclk_obuf_iopad.PULLUP=1'b0;
    defparam apuclk_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD apuclk_obuf_iopad (
            .OE(N__3535),
            .DIN(N__3534),
            .DOUT(N__3533),
            .PACKAGEPIN(apuclk));
    defparam apuclk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam apuclk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO apuclk_obuf_preio (
            .PADOEN(N__3535),
            .PADOUT(N__3534),
            .PADIN(N__3533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3015),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol4_obuf_iopad (
            .OE(N__3526),
            .DIN(N__3525),
            .DOUT(N__3524),
            .PACKAGEPIN(lcol4));
    defparam lcol4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol4_obuf_preio (
            .PADOEN(N__3526),
            .PADOUT(N__3525),
            .PADIN(N__3524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3398),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led2_obuf_iopad (
            .OE(N__3517),
            .DIN(N__3516),
            .DOUT(N__3515),
            .PACKAGEPIN(led2));
    defparam led2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led2_obuf_preio (
            .PADOEN(N__3517),
            .PADOUT(N__3516),
            .PADIN(N__3515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3394),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led4_obuft_iopad (
            .OE(N__3508),
            .DIN(N__3507),
            .DOUT(N__3506),
            .PACKAGEPIN(led4));
    defparam led4_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led4_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led4_obuft_preio (
            .PADOEN(N__3508),
            .PADOUT(N__3507),
            .PADIN(N__3506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led6_obuft_iopad (
            .OE(N__3499),
            .DIN(N__3498),
            .DOUT(N__3497),
            .PACKAGEPIN(led6));
    defparam led6_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led6_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led6_obuft_preio (
            .PADOEN(N__3499),
            .PADOUT(N__3498),
            .PADIN(N__3497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.diveight.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.diveight.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.diveight.io_0_iopad  (
            .OE(N__3490),
            .DIN(N__3489),
            .DOUT(N__3488),
            .PACKAGEPIN(cpuclk));
    defparam \arse.diveight.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.diveight.io_0_preio  (
            .PADOEN(N__3490),
            .PADOUT(N__3489),
            .PADIN(N__3488),
            .CLOCKENABLE(),
            .DOUT1(N__2958),
            .OUTPUTENABLE(N__3390),
            .DIN0(),
            .DOUT0(N__1746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__2949));
    defparam apureset_obuf_iopad.PULLUP=1'b0;
    defparam apureset_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD apureset_obuf_iopad (
            .OE(N__3481),
            .DIN(N__3480),
            .DOUT(N__3479),
            .PACKAGEPIN(apureset));
    defparam apureset_obuf_preio.NEG_TRIGGER=1'b0;
    defparam apureset_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO apureset_obuf_preio (
            .PADOEN(N__3481),
            .PADOUT(N__3480),
            .PADIN(N__3479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3268),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD consolereset_ibuf_iopad (
            .OE(N__3472),
            .DIN(N__3471),
            .DOUT(N__3470),
            .PACKAGEPIN(consolereset));
    defparam consolereset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam consolereset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO consolereset_ibuf_preio (
            .PADOEN(N__3472),
            .PADOUT(N__3471),
            .PADIN(N__3470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(consolereset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol2_obuf_iopad (
            .OE(N__3463),
            .DIN(N__3462),
            .DOUT(N__3461),
            .PACKAGEPIN(lcol2));
    defparam lcol2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol2_obuf_preio (
            .PADOEN(N__3463),
            .PADOUT(N__3462),
            .PADIN(N__3461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led1_obuf_iopad (
            .OE(N__3454),
            .DIN(N__3453),
            .DOUT(N__3452),
            .PACKAGEPIN(led1));
    defparam led1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led1_obuf_preio (
            .PADOEN(N__3454),
            .PADOUT(N__3453),
            .PADIN(N__3452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD apusync_ibuf_iopad (
            .OE(N__3445),
            .DIN(N__3444),
            .DOUT(N__3443),
            .PACKAGEPIN(apusync));
    defparam apusync_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam apusync_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO apusync_ibuf_preio (
            .PADOEN(N__3445),
            .PADOUT(N__3444),
            .PADIN(N__3443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(apusync_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led3_obuft_iopad (
            .OE(N__3436),
            .DIN(N__3435),
            .DOUT(N__3434),
            .PACKAGEPIN(led3));
    defparam led3_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led3_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led3_obuft_preio (
            .PADOEN(N__3436),
            .PADOUT(N__3435),
            .PADIN(N__3434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led5_obuft_iopad (
            .OE(N__3427),
            .DIN(N__3426),
            .DOUT(N__3425),
            .PACKAGEPIN(led5));
    defparam led5_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led5_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led5_obuft_preio (
            .PADOEN(N__3427),
            .PADOUT(N__3426),
            .PADIN(N__3425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led7_obuft_iopad (
            .OE(N__3418),
            .DIN(N__3417),
            .DOUT(N__3416),
            .PACKAGEPIN(led7));
    defparam led7_obuft_preio.NEG_TRIGGER=1'b0;
    defparam led7_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO led7_obuft_preio (
            .PADOEN(N__3418),
            .PADOUT(N__3417),
            .PADIN(N__3416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__798 (
            .O(N__3399),
            .I(N__3395));
    IoInMux I__797 (
            .O(N__3398),
            .I(N__3391));
    LocalMux I__796 (
            .O(N__3395),
            .I(N__3386));
    IoInMux I__795 (
            .O(N__3394),
            .I(N__3383));
    LocalMux I__794 (
            .O(N__3391),
            .I(N__3380));
    IoInMux I__793 (
            .O(N__3390),
            .I(N__3376));
    IoInMux I__792 (
            .O(N__3389),
            .I(N__3373));
    IoSpan4Mux I__791 (
            .O(N__3386),
            .I(N__3367));
    LocalMux I__790 (
            .O(N__3383),
            .I(N__3367));
    IoSpan4Mux I__789 (
            .O(N__3380),
            .I(N__3364));
    IoInMux I__788 (
            .O(N__3379),
            .I(N__3361));
    LocalMux I__787 (
            .O(N__3376),
            .I(N__3358));
    LocalMux I__786 (
            .O(N__3373),
            .I(N__3355));
    InMux I__785 (
            .O(N__3372),
            .I(N__3352));
    IoSpan4Mux I__784 (
            .O(N__3367),
            .I(N__3349));
    IoSpan4Mux I__783 (
            .O(N__3364),
            .I(N__3344));
    LocalMux I__782 (
            .O(N__3361),
            .I(N__3344));
    IoSpan4Mux I__781 (
            .O(N__3358),
            .I(N__3341));
    Span4Mux_s0_h I__780 (
            .O(N__3355),
            .I(N__3338));
    LocalMux I__779 (
            .O(N__3352),
            .I(N__3335));
    IoSpan4Mux I__778 (
            .O(N__3349),
            .I(N__3330));
    IoSpan4Mux I__777 (
            .O(N__3344),
            .I(N__3330));
    Span4Mux_s3_h I__776 (
            .O(N__3341),
            .I(N__3327));
    Span4Mux_h I__775 (
            .O(N__3338),
            .I(N__3322));
    Span4Mux_v I__774 (
            .O(N__3335),
            .I(N__3322));
    Span4Mux_s2_v I__773 (
            .O(N__3330),
            .I(N__3319));
    Sp12to4 I__772 (
            .O(N__3327),
            .I(N__3316));
    Sp12to4 I__771 (
            .O(N__3322),
            .I(N__3313));
    Sp12to4 I__770 (
            .O(N__3319),
            .I(N__3310));
    Span12Mux_h I__769 (
            .O(N__3316),
            .I(N__3305));
    Span12Mux_h I__768 (
            .O(N__3313),
            .I(N__3305));
    Span12Mux_s8_v I__767 (
            .O(N__3310),
            .I(N__3302));
    Odrv12 I__766 (
            .O(N__3305),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__765 (
            .O(N__3302),
            .I(CONSTANT_ONE_NET));
    CEMux I__764 (
            .O(N__3297),
            .I(N__3294));
    LocalMux I__763 (
            .O(N__3294),
            .I(\arse.ddd.N_33_0 ));
    SRMux I__762 (
            .O(N__3291),
            .I(N__3288));
    LocalMux I__761 (
            .O(N__3288),
            .I(N__3285));
    Span4Mux_h I__760 (
            .O(N__3285),
            .I(N__3281));
    InMux I__759 (
            .O(N__3284),
            .I(N__3278));
    Odrv4 I__758 (
            .O(N__3281),
            .I(\arse.seqreset_e_0_RNIQTPZ0Z13 ));
    LocalMux I__757 (
            .O(N__3278),
            .I(\arse.seqreset_e_0_RNIQTPZ0Z13 ));
    CascadeMux I__756 (
            .O(N__3273),
            .I(N__3270));
    InMux I__755 (
            .O(N__3270),
            .I(N__3265));
    InMux I__754 (
            .O(N__3269),
            .I(N__3262));
    IoInMux I__753 (
            .O(N__3268),
            .I(N__3259));
    LocalMux I__752 (
            .O(N__3265),
            .I(N__3256));
    LocalMux I__751 (
            .O(N__3262),
            .I(N__3252));
    LocalMux I__750 (
            .O(N__3259),
            .I(N__3249));
    Span4Mux_v I__749 (
            .O(N__3256),
            .I(N__3246));
    InMux I__748 (
            .O(N__3255),
            .I(N__3243));
    Span4Mux_v I__747 (
            .O(N__3252),
            .I(N__3240));
    Span12Mux_s11_h I__746 (
            .O(N__3249),
            .I(N__3232));
    Sp12to4 I__745 (
            .O(N__3246),
            .I(N__3232));
    LocalMux I__744 (
            .O(N__3243),
            .I(N__3232));
    Span4Mux_h I__743 (
            .O(N__3240),
            .I(N__3229));
    InMux I__742 (
            .O(N__3239),
            .I(N__3226));
    Odrv12 I__741 (
            .O(N__3232),
            .I(apureset_c));
    Odrv4 I__740 (
            .O(N__3229),
            .I(apureset_c));
    LocalMux I__739 (
            .O(N__3226),
            .I(apureset_c));
    InMux I__738 (
            .O(N__3219),
            .I(N__3215));
    InMux I__737 (
            .O(N__3218),
            .I(N__3212));
    LocalMux I__736 (
            .O(N__3215),
            .I(G_73));
    LocalMux I__735 (
            .O(N__3212),
            .I(G_73));
    InMux I__734 (
            .O(N__3207),
            .I(N__3203));
    InMux I__733 (
            .O(N__3206),
            .I(N__3200));
    LocalMux I__732 (
            .O(N__3203),
            .I(N__3194));
    LocalMux I__731 (
            .O(N__3200),
            .I(N__3194));
    InMux I__730 (
            .O(N__3199),
            .I(N__3191));
    Sp12to4 I__729 (
            .O(N__3194),
            .I(N__3186));
    LocalMux I__728 (
            .O(N__3191),
            .I(N__3186));
    Span12Mux_v I__727 (
            .O(N__3186),
            .I(N__3183));
    Span12Mux_h I__726 (
            .O(N__3183),
            .I(N__3180));
    Odrv12 I__725 (
            .O(N__3180),
            .I(apusync_c));
    IoInMux I__724 (
            .O(N__3177),
            .I(N__3174));
    LocalMux I__723 (
            .O(N__3174),
            .I(N__3171));
    IoSpan4Mux I__722 (
            .O(N__3171),
            .I(N__3168));
    Span4Mux_s2_h I__721 (
            .O(N__3168),
            .I(N__3165));
    Span4Mux_h I__720 (
            .O(N__3165),
            .I(N__3161));
    CascadeMux I__719 (
            .O(N__3164),
            .I(N__3158));
    Span4Mux_h I__718 (
            .O(N__3161),
            .I(N__3155));
    InMux I__717 (
            .O(N__3158),
            .I(N__3152));
    Odrv4 I__716 (
            .O(N__3155),
            .I(cpureset_c));
    LocalMux I__715 (
            .O(N__3152),
            .I(cpureset_c));
    InMux I__714 (
            .O(N__3147),
            .I(N__3143));
    CascadeMux I__713 (
            .O(N__3146),
            .I(N__3140));
    LocalMux I__712 (
            .O(N__3143),
            .I(N__3134));
    InMux I__711 (
            .O(N__3140),
            .I(N__3131));
    InMux I__710 (
            .O(N__3139),
            .I(N__3122));
    InMux I__709 (
            .O(N__3138),
            .I(N__3117));
    InMux I__708 (
            .O(N__3137),
            .I(N__3117));
    Span4Mux_v I__707 (
            .O(N__3134),
            .I(N__3114));
    LocalMux I__706 (
            .O(N__3131),
            .I(N__3111));
    InMux I__705 (
            .O(N__3130),
            .I(N__3108));
    InMux I__704 (
            .O(N__3129),
            .I(N__3105));
    InMux I__703 (
            .O(N__3128),
            .I(N__3098));
    InMux I__702 (
            .O(N__3127),
            .I(N__3098));
    InMux I__701 (
            .O(N__3126),
            .I(N__3098));
    InMux I__700 (
            .O(N__3125),
            .I(N__3093));
    LocalMux I__699 (
            .O(N__3122),
            .I(N__3088));
    LocalMux I__698 (
            .O(N__3117),
            .I(N__3088));
    Sp12to4 I__697 (
            .O(N__3114),
            .I(N__3083));
    Span12Mux_s5_v I__696 (
            .O(N__3111),
            .I(N__3083));
    LocalMux I__695 (
            .O(N__3108),
            .I(N__3080));
    LocalMux I__694 (
            .O(N__3105),
            .I(N__3075));
    LocalMux I__693 (
            .O(N__3098),
            .I(N__3075));
    InMux I__692 (
            .O(N__3097),
            .I(N__3069));
    InMux I__691 (
            .O(N__3096),
            .I(N__3069));
    LocalMux I__690 (
            .O(N__3093),
            .I(N__3066));
    Span4Mux_h I__689 (
            .O(N__3088),
            .I(N__3063));
    Span12Mux_h I__688 (
            .O(N__3083),
            .I(N__3060));
    Span4Mux_h I__687 (
            .O(N__3080),
            .I(N__3057));
    Span12Mux_h I__686 (
            .O(N__3075),
            .I(N__3054));
    InMux I__685 (
            .O(N__3074),
            .I(N__3051));
    LocalMux I__684 (
            .O(N__3069),
            .I(\arse.seqresetZ0 ));
    Odrv4 I__683 (
            .O(N__3066),
            .I(\arse.seqresetZ0 ));
    Odrv4 I__682 (
            .O(N__3063),
            .I(\arse.seqresetZ0 ));
    Odrv12 I__681 (
            .O(N__3060),
            .I(\arse.seqresetZ0 ));
    Odrv4 I__680 (
            .O(N__3057),
            .I(\arse.seqresetZ0 ));
    Odrv12 I__679 (
            .O(N__3054),
            .I(\arse.seqresetZ0 ));
    LocalMux I__678 (
            .O(N__3051),
            .I(\arse.seqresetZ0 ));
    InMux I__677 (
            .O(N__3036),
            .I(N__3033));
    LocalMux I__676 (
            .O(N__3033),
            .I(G_74));
    InMux I__675 (
            .O(N__3030),
            .I(N__3027));
    LocalMux I__674 (
            .O(N__3027),
            .I(N__3024));
    Span12Mux_h I__673 (
            .O(N__3024),
            .I(N__3021));
    Odrv12 I__672 (
            .O(N__3021),
            .I(\arse.divseven.io_0_D_IN_0 ));
    CascadeMux I__671 (
            .O(N__3018),
            .I(G_74_cascade_));
    IoInMux I__670 (
            .O(N__3015),
            .I(N__3012));
    LocalMux I__669 (
            .O(N__3012),
            .I(N__3009));
    IoSpan4Mux I__668 (
            .O(N__3009),
            .I(N__3006));
    Span4Mux_s3_h I__667 (
            .O(N__3006),
            .I(N__3003));
    Span4Mux_v I__666 (
            .O(N__3003),
            .I(N__3000));
    Sp12to4 I__665 (
            .O(N__3000),
            .I(N__2997));
    Odrv12 I__664 (
            .O(N__2997),
            .I(arse_un1_apuclk_i));
    InMux I__663 (
            .O(N__2994),
            .I(N__2991));
    LocalMux I__662 (
            .O(N__2991),
            .I(N__2988));
    Span4Mux_v I__661 (
            .O(N__2988),
            .I(N__2985));
    Sp12to4 I__660 (
            .O(N__2985),
            .I(N__2982));
    Span12Mux_s5_h I__659 (
            .O(N__2982),
            .I(N__2978));
    InMux I__658 (
            .O(N__2981),
            .I(N__2974));
    Span12Mux_h I__657 (
            .O(N__2978),
            .I(N__2971));
    InMux I__656 (
            .O(N__2977),
            .I(N__2968));
    LocalMux I__655 (
            .O(N__2974),
            .I(N__2965));
    Odrv12 I__654 (
            .O(N__2971),
            .I(\arse.diveight.counterZ0Z_2 ));
    LocalMux I__653 (
            .O(N__2968),
            .I(\arse.diveight.counterZ0Z_2 ));
    Odrv4 I__652 (
            .O(N__2965),
            .I(\arse.diveight.counterZ0Z_2 ));
    IoInMux I__651 (
            .O(N__2958),
            .I(N__2955));
    LocalMux I__650 (
            .O(N__2955),
            .I(N__2952));
    Odrv4 I__649 (
            .O(N__2952),
            .I(\arse.diveight.doutZ0Z_1 ));
    ClkMux I__648 (
            .O(N__2949),
            .I(N__2898));
    ClkMux I__647 (
            .O(N__2948),
            .I(N__2898));
    ClkMux I__646 (
            .O(N__2947),
            .I(N__2898));
    ClkMux I__645 (
            .O(N__2946),
            .I(N__2898));
    ClkMux I__644 (
            .O(N__2945),
            .I(N__2898));
    ClkMux I__643 (
            .O(N__2944),
            .I(N__2898));
    ClkMux I__642 (
            .O(N__2943),
            .I(N__2898));
    ClkMux I__641 (
            .O(N__2942),
            .I(N__2898));
    ClkMux I__640 (
            .O(N__2941),
            .I(N__2898));
    ClkMux I__639 (
            .O(N__2940),
            .I(N__2898));
    ClkMux I__638 (
            .O(N__2939),
            .I(N__2898));
    ClkMux I__637 (
            .O(N__2938),
            .I(N__2898));
    ClkMux I__636 (
            .O(N__2937),
            .I(N__2898));
    ClkMux I__635 (
            .O(N__2936),
            .I(N__2898));
    ClkMux I__634 (
            .O(N__2935),
            .I(N__2898));
    ClkMux I__633 (
            .O(N__2934),
            .I(N__2898));
    ClkMux I__632 (
            .O(N__2933),
            .I(N__2898));
    GlobalMux I__631 (
            .O(N__2898),
            .I(N__2895));
    gio2CtrlBuf I__630 (
            .O(N__2895),
            .I(PLLOUTCORE_0_g));
    SRMux I__629 (
            .O(N__2892),
            .I(N__2889));
    LocalMux I__628 (
            .O(N__2889),
            .I(N__2884));
    SRMux I__627 (
            .O(N__2888),
            .I(N__2881));
    SRMux I__626 (
            .O(N__2887),
            .I(N__2876));
    Span4Mux_s3_h I__625 (
            .O(N__2884),
            .I(N__2873));
    LocalMux I__624 (
            .O(N__2881),
            .I(N__2870));
    SRMux I__623 (
            .O(N__2880),
            .I(N__2867));
    SRMux I__622 (
            .O(N__2879),
            .I(N__2863));
    LocalMux I__621 (
            .O(N__2876),
            .I(N__2860));
    Sp12to4 I__620 (
            .O(N__2873),
            .I(N__2857));
    Span4Mux_v I__619 (
            .O(N__2870),
            .I(N__2852));
    LocalMux I__618 (
            .O(N__2867),
            .I(N__2852));
    SRMux I__617 (
            .O(N__2866),
            .I(N__2849));
    LocalMux I__616 (
            .O(N__2863),
            .I(N__2846));
    Span4Mux_s0_v I__615 (
            .O(N__2860),
            .I(N__2843));
    Span12Mux_h I__614 (
            .O(N__2857),
            .I(N__2834));
    Sp12to4 I__613 (
            .O(N__2852),
            .I(N__2834));
    LocalMux I__612 (
            .O(N__2849),
            .I(N__2834));
    Span4Mux_h I__611 (
            .O(N__2846),
            .I(N__2831));
    Span4Mux_h I__610 (
            .O(N__2843),
            .I(N__2828));
    SRMux I__609 (
            .O(N__2842),
            .I(N__2825));
    InMux I__608 (
            .O(N__2841),
            .I(N__2822));
    Odrv12 I__607 (
            .O(N__2834),
            .I(\arse.seqreset_i ));
    Odrv4 I__606 (
            .O(N__2831),
            .I(\arse.seqreset_i ));
    Odrv4 I__605 (
            .O(N__2828),
            .I(\arse.seqreset_i ));
    LocalMux I__604 (
            .O(N__2825),
            .I(\arse.seqreset_i ));
    LocalMux I__603 (
            .O(N__2822),
            .I(\arse.seqreset_i ));
    InMux I__602 (
            .O(N__2811),
            .I(N__2805));
    InMux I__601 (
            .O(N__2810),
            .I(N__2802));
    InMux I__600 (
            .O(N__2809),
            .I(N__2799));
    InMux I__599 (
            .O(N__2808),
            .I(N__2796));
    LocalMux I__598 (
            .O(N__2805),
            .I(\arse.arse.counterZ0Z_2 ));
    LocalMux I__597 (
            .O(N__2802),
            .I(\arse.arse.counterZ0Z_2 ));
    LocalMux I__596 (
            .O(N__2799),
            .I(\arse.arse.counterZ0Z_2 ));
    LocalMux I__595 (
            .O(N__2796),
            .I(\arse.arse.counterZ0Z_2 ));
    CascadeMux I__594 (
            .O(N__2787),
            .I(N__2784));
    InMux I__593 (
            .O(N__2784),
            .I(N__2781));
    LocalMux I__592 (
            .O(N__2781),
            .I(\arse.arse.un16_counter_cry_1_THRU_CO ));
    InMux I__591 (
            .O(N__2778),
            .I(\arse.arse.un16_counter_cry_1 ));
    CascadeMux I__590 (
            .O(N__2775),
            .I(N__2772));
    InMux I__589 (
            .O(N__2772),
            .I(N__2769));
    LocalMux I__588 (
            .O(N__2769),
            .I(\arse.arse.un16_counter_cry_2_THRU_CO ));
    InMux I__587 (
            .O(N__2766),
            .I(\arse.arse.un16_counter_cry_2 ));
    InMux I__586 (
            .O(N__2763),
            .I(\arse.arse.un16_counter_cry_3 ));
    InMux I__585 (
            .O(N__2760),
            .I(N__2756));
    InMux I__584 (
            .O(N__2759),
            .I(N__2753));
    LocalMux I__583 (
            .O(N__2756),
            .I(\arse.arse.counterZ0Z_4 ));
    LocalMux I__582 (
            .O(N__2753),
            .I(\arse.arse.counterZ0Z_4 ));
    InMux I__581 (
            .O(N__2748),
            .I(N__2743));
    InMux I__580 (
            .O(N__2747),
            .I(N__2740));
    InMux I__579 (
            .O(N__2746),
            .I(N__2737));
    LocalMux I__578 (
            .O(N__2743),
            .I(\arse.arse.counterZ0Z_3 ));
    LocalMux I__577 (
            .O(N__2740),
            .I(\arse.arse.counterZ0Z_3 ));
    LocalMux I__576 (
            .O(N__2737),
            .I(\arse.arse.counterZ0Z_3 ));
    CascadeMux I__575 (
            .O(N__2730),
            .I(\arse.G_2_0_cascade_ ));
    InMux I__574 (
            .O(N__2727),
            .I(N__2721));
    InMux I__573 (
            .O(N__2726),
            .I(N__2721));
    LocalMux I__572 (
            .O(N__2721),
            .I(N__2718));
    Span4Mux_v I__571 (
            .O(N__2718),
            .I(N__2709));
    InMux I__570 (
            .O(N__2717),
            .I(N__2706));
    InMux I__569 (
            .O(N__2716),
            .I(N__2703));
    InMux I__568 (
            .O(N__2715),
            .I(N__2700));
    InMux I__567 (
            .O(N__2714),
            .I(N__2693));
    InMux I__566 (
            .O(N__2713),
            .I(N__2693));
    InMux I__565 (
            .O(N__2712),
            .I(N__2693));
    Odrv4 I__564 (
            .O(N__2709),
            .I(\arse.un1_counterlto4_0 ));
    LocalMux I__563 (
            .O(N__2706),
            .I(\arse.un1_counterlto4_0 ));
    LocalMux I__562 (
            .O(N__2703),
            .I(\arse.un1_counterlto4_0 ));
    LocalMux I__561 (
            .O(N__2700),
            .I(\arse.un1_counterlto4_0 ));
    LocalMux I__560 (
            .O(N__2693),
            .I(\arse.un1_counterlto4_0 ));
    CascadeMux I__559 (
            .O(N__2682),
            .I(N__2679));
    InMux I__558 (
            .O(N__2679),
            .I(N__2672));
    InMux I__557 (
            .O(N__2678),
            .I(N__2663));
    InMux I__556 (
            .O(N__2677),
            .I(N__2663));
    InMux I__555 (
            .O(N__2676),
            .I(N__2663));
    InMux I__554 (
            .O(N__2675),
            .I(N__2660));
    LocalMux I__553 (
            .O(N__2672),
            .I(N__2657));
    InMux I__552 (
            .O(N__2671),
            .I(N__2652));
    InMux I__551 (
            .O(N__2670),
            .I(N__2652));
    LocalMux I__550 (
            .O(N__2663),
            .I(N__2649));
    LocalMux I__549 (
            .O(N__2660),
            .I(\arse.un1_counterlt4 ));
    Odrv4 I__548 (
            .O(N__2657),
            .I(\arse.un1_counterlt4 ));
    LocalMux I__547 (
            .O(N__2652),
            .I(\arse.un1_counterlt4 ));
    Odrv4 I__546 (
            .O(N__2649),
            .I(\arse.un1_counterlt4 ));
    CascadeMux I__545 (
            .O(N__2640),
            .I(N__2636));
    CascadeMux I__544 (
            .O(N__2639),
            .I(N__2633));
    InMux I__543 (
            .O(N__2636),
            .I(N__2625));
    InMux I__542 (
            .O(N__2633),
            .I(N__2625));
    InMux I__541 (
            .O(N__2632),
            .I(N__2625));
    LocalMux I__540 (
            .O(N__2625),
            .I(\arse.clock_out_i ));
    InMux I__539 (
            .O(N__2622),
            .I(N__2619));
    LocalMux I__538 (
            .O(N__2619),
            .I(\arse.ddd.Q_esr_RNOZ0Z_0 ));
    InMux I__537 (
            .O(N__2616),
            .I(N__2613));
    LocalMux I__536 (
            .O(N__2613),
            .I(N__2610));
    Span12Mux_v I__535 (
            .O(N__2610),
            .I(N__2607));
    Span12Mux_v I__534 (
            .O(N__2607),
            .I(N__2604));
    Odrv12 I__533 (
            .O(N__2604),
            .I(consolereset_c));
    CascadeMux I__532 (
            .O(N__2601),
            .I(\debounceconsolereset.out_cnv_4_cascade_ ));
    CascadeMux I__531 (
            .O(N__2598),
            .I(N__2592));
    InMux I__530 (
            .O(N__2597),
            .I(N__2583));
    InMux I__529 (
            .O(N__2596),
            .I(N__2583));
    InMux I__528 (
            .O(N__2595),
            .I(N__2580));
    InMux I__527 (
            .O(N__2592),
            .I(N__2575));
    InMux I__526 (
            .O(N__2591),
            .I(N__2575));
    InMux I__525 (
            .O(N__2590),
            .I(N__2568));
    InMux I__524 (
            .O(N__2589),
            .I(N__2568));
    InMux I__523 (
            .O(N__2588),
            .I(N__2568));
    LocalMux I__522 (
            .O(N__2583),
            .I(clock_out_RNIR6ER));
    LocalMux I__521 (
            .O(N__2580),
            .I(clock_out_RNIR6ER));
    LocalMux I__520 (
            .O(N__2575),
            .I(clock_out_RNIR6ER));
    LocalMux I__519 (
            .O(N__2568),
            .I(clock_out_RNIR6ER));
    CascadeMux I__518 (
            .O(N__2559),
            .I(N__2556));
    InMux I__517 (
            .O(N__2556),
            .I(N__2547));
    InMux I__516 (
            .O(N__2555),
            .I(N__2542));
    InMux I__515 (
            .O(N__2554),
            .I(N__2542));
    InMux I__514 (
            .O(N__2553),
            .I(N__2533));
    InMux I__513 (
            .O(N__2552),
            .I(N__2533));
    InMux I__512 (
            .O(N__2551),
            .I(N__2533));
    InMux I__511 (
            .O(N__2550),
            .I(N__2533));
    LocalMux I__510 (
            .O(N__2547),
            .I(\debounceconsolereset.counter_RNI4RTH1Z0Z_6 ));
    LocalMux I__509 (
            .O(N__2542),
            .I(\debounceconsolereset.counter_RNI4RTH1Z0Z_6 ));
    LocalMux I__508 (
            .O(N__2533),
            .I(\debounceconsolereset.counter_RNI4RTH1Z0Z_6 ));
    InMux I__507 (
            .O(N__2526),
            .I(N__2522));
    CascadeMux I__506 (
            .O(N__2525),
            .I(N__2517));
    LocalMux I__505 (
            .O(N__2522),
            .I(N__2514));
    InMux I__504 (
            .O(N__2521),
            .I(N__2509));
    InMux I__503 (
            .O(N__2520),
            .I(N__2509));
    InMux I__502 (
            .O(N__2517),
            .I(N__2506));
    Odrv4 I__501 (
            .O(N__2514),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    LocalMux I__500 (
            .O(N__2509),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    LocalMux I__499 (
            .O(N__2506),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    CascadeMux I__498 (
            .O(N__2499),
            .I(N__2495));
    CascadeMux I__497 (
            .O(N__2498),
            .I(N__2492));
    InMux I__496 (
            .O(N__2495),
            .I(N__2486));
    InMux I__495 (
            .O(N__2492),
            .I(N__2486));
    InMux I__494 (
            .O(N__2491),
            .I(N__2483));
    LocalMux I__493 (
            .O(N__2486),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    LocalMux I__492 (
            .O(N__2483),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    InMux I__491 (
            .O(N__2478),
            .I(N__2475));
    LocalMux I__490 (
            .O(N__2475),
            .I(N__2466));
    ClkMux I__489 (
            .O(N__2474),
            .I(N__2451));
    ClkMux I__488 (
            .O(N__2473),
            .I(N__2451));
    ClkMux I__487 (
            .O(N__2472),
            .I(N__2451));
    ClkMux I__486 (
            .O(N__2471),
            .I(N__2451));
    ClkMux I__485 (
            .O(N__2470),
            .I(N__2451));
    ClkMux I__484 (
            .O(N__2469),
            .I(N__2451));
    Glb2LocalMux I__483 (
            .O(N__2466),
            .I(N__2451));
    GlobalMux I__482 (
            .O(N__2451),
            .I(N__2448));
    gio2CtrlBuf I__481 (
            .O(N__2448),
            .I(PACKAGEPIN_0_c_g));
    IoInMux I__480 (
            .O(N__2445),
            .I(N__2442));
    LocalMux I__479 (
            .O(N__2442),
            .I(N__2439));
    IoSpan4Mux I__478 (
            .O(N__2439),
            .I(N__2436));
    Odrv4 I__477 (
            .O(N__2436),
            .I(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO));
    InMux I__476 (
            .O(N__2433),
            .I(N__2427));
    InMux I__475 (
            .O(N__2432),
            .I(N__2424));
    InMux I__474 (
            .O(N__2431),
            .I(N__2421));
    InMux I__473 (
            .O(N__2430),
            .I(N__2418));
    LocalMux I__472 (
            .O(N__2427),
            .I(\arse.arse.counterZ0Z_0 ));
    LocalMux I__471 (
            .O(N__2424),
            .I(\arse.arse.counterZ0Z_0 ));
    LocalMux I__470 (
            .O(N__2421),
            .I(\arse.arse.counterZ0Z_0 ));
    LocalMux I__469 (
            .O(N__2418),
            .I(\arse.arse.counterZ0Z_0 ));
    CascadeMux I__468 (
            .O(N__2409),
            .I(N__2405));
    CascadeMux I__467 (
            .O(N__2408),
            .I(N__2402));
    InMux I__466 (
            .O(N__2405),
            .I(N__2398));
    InMux I__465 (
            .O(N__2402),
            .I(N__2395));
    InMux I__464 (
            .O(N__2401),
            .I(N__2392));
    LocalMux I__463 (
            .O(N__2398),
            .I(\arse.arse.counterZ0Z_1 ));
    LocalMux I__462 (
            .O(N__2395),
            .I(\arse.arse.counterZ0Z_1 ));
    LocalMux I__461 (
            .O(N__2392),
            .I(\arse.arse.counterZ0Z_1 ));
    InMux I__460 (
            .O(N__2385),
            .I(N__2382));
    LocalMux I__459 (
            .O(N__2382),
            .I(\debounceconsolereset.un3_counter_cry_2_THRU_CO ));
    InMux I__458 (
            .O(N__2379),
            .I(\debounceconsolereset.un3_counter_cry_2 ));
    InMux I__457 (
            .O(N__2376),
            .I(N__2370));
    InMux I__456 (
            .O(N__2375),
            .I(N__2363));
    InMux I__455 (
            .O(N__2374),
            .I(N__2363));
    InMux I__454 (
            .O(N__2373),
            .I(N__2363));
    LocalMux I__453 (
            .O(N__2370),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    LocalMux I__452 (
            .O(N__2363),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    InMux I__451 (
            .O(N__2358),
            .I(N__2355));
    LocalMux I__450 (
            .O(N__2355),
            .I(\debounceconsolereset.un3_counter_cry_3_THRU_CO ));
    InMux I__449 (
            .O(N__2352),
            .I(\debounceconsolereset.un3_counter_cry_3 ));
    InMux I__448 (
            .O(N__2349),
            .I(\debounceconsolereset.un3_counter_cry_4 ));
    InMux I__447 (
            .O(N__2346),
            .I(\debounceconsolereset.un3_counter_cry_5 ));
    CascadeMux I__446 (
            .O(N__2343),
            .I(clock_out_RNIR6ER_cascade_));
    InMux I__445 (
            .O(N__2340),
            .I(N__2337));
    LocalMux I__444 (
            .O(N__2337),
            .I(\debounceconsolereset.un1_counterlt6 ));
    InMux I__443 (
            .O(N__2334),
            .I(N__2330));
    InMux I__442 (
            .O(N__2333),
            .I(N__2327));
    LocalMux I__441 (
            .O(N__2330),
            .I(N__2322));
    LocalMux I__440 (
            .O(N__2327),
            .I(N__2319));
    InMux I__439 (
            .O(N__2326),
            .I(N__2315));
    CEMux I__438 (
            .O(N__2325),
            .I(N__2312));
    Span4Mux_v I__437 (
            .O(N__2322),
            .I(N__2304));
    Span4Mux_v I__436 (
            .O(N__2319),
            .I(N__2301));
    IoInMux I__435 (
            .O(N__2318),
            .I(N__2298));
    LocalMux I__434 (
            .O(N__2315),
            .I(N__2295));
    LocalMux I__433 (
            .O(N__2312),
            .I(N__2292));
    InMux I__432 (
            .O(N__2311),
            .I(N__2285));
    InMux I__431 (
            .O(N__2310),
            .I(N__2285));
    InMux I__430 (
            .O(N__2309),
            .I(N__2285));
    InMux I__429 (
            .O(N__2308),
            .I(N__2280));
    InMux I__428 (
            .O(N__2307),
            .I(N__2280));
    Span4Mux_h I__427 (
            .O(N__2304),
            .I(N__2275));
    Span4Mux_h I__426 (
            .O(N__2301),
            .I(N__2275));
    LocalMux I__425 (
            .O(N__2298),
            .I(N__2272));
    Span4Mux_v I__424 (
            .O(N__2295),
            .I(N__2269));
    Span4Mux_v I__423 (
            .O(N__2292),
            .I(N__2262));
    LocalMux I__422 (
            .O(N__2285),
            .I(N__2262));
    LocalMux I__421 (
            .O(N__2280),
            .I(N__2262));
    Span4Mux_h I__420 (
            .O(N__2275),
            .I(N__2257));
    Span4Mux_s2_v I__419 (
            .O(N__2272),
            .I(N__2257));
    Sp12to4 I__418 (
            .O(N__2269),
            .I(N__2254));
    Span4Mux_v I__417 (
            .O(N__2262),
            .I(N__2251));
    Span4Mux_h I__416 (
            .O(N__2257),
            .I(N__2248));
    Span12Mux_h I__415 (
            .O(N__2254),
            .I(N__2245));
    Sp12to4 I__414 (
            .O(N__2251),
            .I(N__2242));
    Span4Mux_h I__413 (
            .O(N__2248),
            .I(N__2239));
    Span12Mux_h I__412 (
            .O(N__2245),
            .I(N__2236));
    Span12Mux_h I__411 (
            .O(N__2242),
            .I(N__2233));
    Sp12to4 I__410 (
            .O(N__2239),
            .I(N__2230));
    Span12Mux_v I__409 (
            .O(N__2236),
            .I(N__2227));
    Span12Mux_h I__408 (
            .O(N__2233),
            .I(N__2224));
    Span12Mux_v I__407 (
            .O(N__2230),
            .I(N__2221));
    Span12Mux_v I__406 (
            .O(N__2227),
            .I(N__2218));
    Span12Mux_v I__405 (
            .O(N__2224),
            .I(N__2215));
    Span12Mux_v I__404 (
            .O(N__2221),
            .I(N__2212));
    Odrv12 I__403 (
            .O(N__2218),
            .I(masterreset_c));
    Odrv12 I__402 (
            .O(N__2215),
            .I(masterreset_c));
    Odrv12 I__401 (
            .O(N__2212),
            .I(masterreset_c));
    InMux I__400 (
            .O(N__2205),
            .I(N__2186));
    InMux I__399 (
            .O(N__2204),
            .I(N__2177));
    InMux I__398 (
            .O(N__2203),
            .I(N__2177));
    InMux I__397 (
            .O(N__2202),
            .I(N__2177));
    InMux I__396 (
            .O(N__2201),
            .I(N__2177));
    InMux I__395 (
            .O(N__2200),
            .I(N__2170));
    InMux I__394 (
            .O(N__2199),
            .I(N__2170));
    InMux I__393 (
            .O(N__2198),
            .I(N__2170));
    InMux I__392 (
            .O(N__2197),
            .I(N__2165));
    InMux I__391 (
            .O(N__2196),
            .I(N__2165));
    InMux I__390 (
            .O(N__2195),
            .I(N__2158));
    InMux I__389 (
            .O(N__2194),
            .I(N__2158));
    InMux I__388 (
            .O(N__2193),
            .I(N__2158));
    InMux I__387 (
            .O(N__2192),
            .I(N__2151));
    InMux I__386 (
            .O(N__2191),
            .I(N__2151));
    InMux I__385 (
            .O(N__2190),
            .I(N__2151));
    InMux I__384 (
            .O(N__2189),
            .I(N__2148));
    LocalMux I__383 (
            .O(N__2186),
            .I(\arses.counter8 ));
    LocalMux I__382 (
            .O(N__2177),
            .I(\arses.counter8 ));
    LocalMux I__381 (
            .O(N__2170),
            .I(\arses.counter8 ));
    LocalMux I__380 (
            .O(N__2165),
            .I(\arses.counter8 ));
    LocalMux I__379 (
            .O(N__2158),
            .I(\arses.counter8 ));
    LocalMux I__378 (
            .O(N__2151),
            .I(\arses.counter8 ));
    LocalMux I__377 (
            .O(N__2148),
            .I(\arses.counter8 ));
    InMux I__376 (
            .O(N__2133),
            .I(N__2129));
    InMux I__375 (
            .O(N__2132),
            .I(N__2126));
    LocalMux I__374 (
            .O(N__2129),
            .I(\arses.clock_out_i ));
    LocalMux I__373 (
            .O(N__2126),
            .I(\arses.clock_out_i ));
    CascadeMux I__372 (
            .O(N__2121),
            .I(N__2118));
    InMux I__371 (
            .O(N__2118),
            .I(N__2115));
    LocalMux I__370 (
            .O(N__2115),
            .I(\debounceconsolereset.un3_counter_cry_4_THRU_CO ));
    InMux I__369 (
            .O(N__2112),
            .I(N__2104));
    InMux I__368 (
            .O(N__2111),
            .I(N__2104));
    InMux I__367 (
            .O(N__2110),
            .I(N__2099));
    InMux I__366 (
            .O(N__2109),
            .I(N__2099));
    LocalMux I__365 (
            .O(N__2104),
            .I(\debounceconsolereset.counterZ0Z_5 ));
    LocalMux I__364 (
            .O(N__2099),
            .I(\debounceconsolereset.counterZ0Z_5 ));
    InMux I__363 (
            .O(N__2094),
            .I(N__2091));
    LocalMux I__362 (
            .O(N__2091),
            .I(N__2088));
    Odrv4 I__361 (
            .O(N__2088),
            .I(\debounceconsolereset.out_cnv_3 ));
    InMux I__360 (
            .O(N__2085),
            .I(N__2080));
    InMux I__359 (
            .O(N__2084),
            .I(N__2077));
    InMux I__358 (
            .O(N__2083),
            .I(N__2074));
    LocalMux I__357 (
            .O(N__2080),
            .I(\debounceconsolereset.counterZ0Z_6 ));
    LocalMux I__356 (
            .O(N__2077),
            .I(\debounceconsolereset.counterZ0Z_6 ));
    LocalMux I__355 (
            .O(N__2074),
            .I(\debounceconsolereset.counterZ0Z_6 ));
    InMux I__354 (
            .O(N__2067),
            .I(N__2063));
    InMux I__353 (
            .O(N__2066),
            .I(N__2060));
    LocalMux I__352 (
            .O(N__2063),
            .I(\arses.counterZ0Z_14 ));
    LocalMux I__351 (
            .O(N__2060),
            .I(\arses.counterZ0Z_14 ));
    InMux I__350 (
            .O(N__2055),
            .I(N__2051));
    InMux I__349 (
            .O(N__2054),
            .I(N__2048));
    LocalMux I__348 (
            .O(N__2051),
            .I(\arses.counterZ0Z_13 ));
    LocalMux I__347 (
            .O(N__2048),
            .I(\arses.counterZ0Z_13 ));
    CascadeMux I__346 (
            .O(N__2043),
            .I(\arses.un1_counterlt13_0_cascade_ ));
    InMux I__345 (
            .O(N__2040),
            .I(N__2036));
    InMux I__344 (
            .O(N__2039),
            .I(N__2033));
    LocalMux I__343 (
            .O(N__2036),
            .I(\arses.counterZ0Z_12 ));
    LocalMux I__342 (
            .O(N__2033),
            .I(\arses.counterZ0Z_12 ));
    CascadeMux I__341 (
            .O(N__2028),
            .I(N__2025));
    InMux I__340 (
            .O(N__2025),
            .I(N__2015));
    InMux I__339 (
            .O(N__2024),
            .I(N__2015));
    InMux I__338 (
            .O(N__2023),
            .I(N__2015));
    InMux I__337 (
            .O(N__2022),
            .I(N__2012));
    LocalMux I__336 (
            .O(N__2015),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    LocalMux I__335 (
            .O(N__2012),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    InMux I__334 (
            .O(N__2007),
            .I(N__2004));
    LocalMux I__333 (
            .O(N__2004),
            .I(\debounceconsolereset.un3_counter_cry_1_THRU_CO ));
    InMux I__332 (
            .O(N__2001),
            .I(\debounceconsolereset.un3_counter_cry_1 ));
    CascadeMux I__331 (
            .O(N__1998),
            .I(N__1993));
    CascadeMux I__330 (
            .O(N__1997),
            .I(N__1990));
    InMux I__329 (
            .O(N__1996),
            .I(N__1986));
    InMux I__328 (
            .O(N__1993),
            .I(N__1979));
    InMux I__327 (
            .O(N__1990),
            .I(N__1979));
    InMux I__326 (
            .O(N__1989),
            .I(N__1979));
    LocalMux I__325 (
            .O(N__1986),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    LocalMux I__324 (
            .O(N__1979),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    CascadeMux I__323 (
            .O(N__1974),
            .I(N__1971));
    InMux I__322 (
            .O(N__1971),
            .I(N__1965));
    InMux I__321 (
            .O(N__1970),
            .I(N__1965));
    LocalMux I__320 (
            .O(N__1965),
            .I(\arse.diveight.counterZ0Z_1 ));
    CascadeMux I__319 (
            .O(N__1962),
            .I(N__1958));
    InMux I__318 (
            .O(N__1961),
            .I(N__1954));
    InMux I__317 (
            .O(N__1958),
            .I(N__1949));
    InMux I__316 (
            .O(N__1957),
            .I(N__1949));
    LocalMux I__315 (
            .O(N__1954),
            .I(\arse.diveight.counterZ0Z_0 ));
    LocalMux I__314 (
            .O(N__1949),
            .I(\arse.diveight.counterZ0Z_0 ));
    InMux I__313 (
            .O(N__1944),
            .I(N__1940));
    InMux I__312 (
            .O(N__1943),
            .I(N__1937));
    LocalMux I__311 (
            .O(N__1940),
            .I(\arses.counterZ0Z_3 ));
    LocalMux I__310 (
            .O(N__1937),
            .I(\arses.counterZ0Z_3 ));
    InMux I__309 (
            .O(N__1932),
            .I(N__1928));
    InMux I__308 (
            .O(N__1931),
            .I(N__1925));
    LocalMux I__307 (
            .O(N__1928),
            .I(\arses.counterZ0Z_2 ));
    LocalMux I__306 (
            .O(N__1925),
            .I(\arses.counterZ0Z_2 ));
    InMux I__305 (
            .O(N__1920),
            .I(N__1916));
    InMux I__304 (
            .O(N__1919),
            .I(N__1913));
    LocalMux I__303 (
            .O(N__1916),
            .I(N__1910));
    LocalMux I__302 (
            .O(N__1913),
            .I(\arses.counterZ0Z_4 ));
    Odrv4 I__301 (
            .O(N__1910),
            .I(\arses.counterZ0Z_4 ));
    CascadeMux I__300 (
            .O(N__1905),
            .I(\arses.un1_counterlto4_2_cascade_ ));
    InMux I__299 (
            .O(N__1902),
            .I(N__1899));
    LocalMux I__298 (
            .O(N__1899),
            .I(\arses.un1_counterlto8_2 ));
    InMux I__297 (
            .O(N__1896),
            .I(N__1893));
    LocalMux I__296 (
            .O(N__1893),
            .I(N__1887));
    InMux I__295 (
            .O(N__1892),
            .I(N__1880));
    InMux I__294 (
            .O(N__1891),
            .I(N__1880));
    InMux I__293 (
            .O(N__1890),
            .I(N__1880));
    Odrv4 I__292 (
            .O(N__1887),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__291 (
            .O(N__1880),
            .I(\arses.counterZ0Z_0 ));
    CascadeMux I__290 (
            .O(N__1875),
            .I(N__1871));
    CascadeMux I__289 (
            .O(N__1874),
            .I(N__1868));
    InMux I__288 (
            .O(N__1871),
            .I(N__1864));
    InMux I__287 (
            .O(N__1868),
            .I(N__1859));
    InMux I__286 (
            .O(N__1867),
            .I(N__1859));
    LocalMux I__285 (
            .O(N__1864),
            .I(\arses.counterZ0Z_1 ));
    LocalMux I__284 (
            .O(N__1859),
            .I(\arses.counterZ0Z_1 ));
    SRMux I__283 (
            .O(N__1854),
            .I(N__1849));
    SRMux I__282 (
            .O(N__1853),
            .I(N__1846));
    SRMux I__281 (
            .O(N__1852),
            .I(N__1843));
    LocalMux I__280 (
            .O(N__1849),
            .I(N__1840));
    LocalMux I__279 (
            .O(N__1846),
            .I(N__1835));
    LocalMux I__278 (
            .O(N__1843),
            .I(N__1835));
    Span4Mux_v I__277 (
            .O(N__1840),
            .I(N__1832));
    Odrv4 I__276 (
            .O(N__1835),
            .I(masterreset_c_i));
    Odrv4 I__275 (
            .O(N__1832),
            .I(masterreset_c_i));
    InMux I__274 (
            .O(N__1827),
            .I(N__1823));
    InMux I__273 (
            .O(N__1826),
            .I(N__1820));
    LocalMux I__272 (
            .O(N__1823),
            .I(\arses.counterZ0Z_10 ));
    LocalMux I__271 (
            .O(N__1820),
            .I(\arses.counterZ0Z_10 ));
    InMux I__270 (
            .O(N__1815),
            .I(N__1812));
    LocalMux I__269 (
            .O(N__1812),
            .I(\arses.un1_counterlt11 ));
    CascadeMux I__268 (
            .O(N__1809),
            .I(N__1805));
    InMux I__267 (
            .O(N__1808),
            .I(N__1802));
    InMux I__266 (
            .O(N__1805),
            .I(N__1799));
    LocalMux I__265 (
            .O(N__1802),
            .I(\arses.counterZ0Z_11 ));
    LocalMux I__264 (
            .O(N__1799),
            .I(\arses.counterZ0Z_11 ));
    InMux I__263 (
            .O(N__1794),
            .I(N__1790));
    InMux I__262 (
            .O(N__1793),
            .I(N__1787));
    LocalMux I__261 (
            .O(N__1790),
            .I(\arses.counterZ0Z_9 ));
    LocalMux I__260 (
            .O(N__1787),
            .I(\arses.counterZ0Z_9 ));
    CascadeMux I__259 (
            .O(N__1782),
            .I(N__1778));
    InMux I__258 (
            .O(N__1781),
            .I(N__1775));
    InMux I__257 (
            .O(N__1778),
            .I(N__1772));
    LocalMux I__256 (
            .O(N__1775),
            .I(\arses.counterZ0Z_8 ));
    LocalMux I__255 (
            .O(N__1772),
            .I(\arses.counterZ0Z_8 ));
    InMux I__254 (
            .O(N__1767),
            .I(\arses.un2_counter_cry_7 ));
    InMux I__253 (
            .O(N__1764),
            .I(bfn_9_5_0_));
    InMux I__252 (
            .O(N__1761),
            .I(\arses.un2_counter_cry_9 ));
    InMux I__251 (
            .O(N__1758),
            .I(\arses.un2_counter_cry_10 ));
    InMux I__250 (
            .O(N__1755),
            .I(\arses.un2_counter_cry_11 ));
    InMux I__249 (
            .O(N__1752),
            .I(\arses.un2_counter_cry_12 ));
    InMux I__248 (
            .O(N__1749),
            .I(\arses.un2_counter_cry_13 ));
    IoInMux I__247 (
            .O(N__1746),
            .I(N__1743));
    LocalMux I__246 (
            .O(N__1743),
            .I(N__1740));
    Span4Mux_s1_h I__245 (
            .O(N__1740),
            .I(N__1737));
    Span4Mux_v I__244 (
            .O(N__1737),
            .I(N__1734));
    Sp12to4 I__243 (
            .O(N__1734),
            .I(N__1731));
    Span12Mux_h I__242 (
            .O(N__1731),
            .I(N__1728));
    Odrv12 I__241 (
            .O(N__1728),
            .I(\arse.diveight.doutZ0Z_0 ));
    InMux I__240 (
            .O(N__1725),
            .I(N__1722));
    LocalMux I__239 (
            .O(N__1722),
            .I(N__1717));
    InMux I__238 (
            .O(N__1721),
            .I(N__1712));
    InMux I__237 (
            .O(N__1720),
            .I(N__1712));
    Odrv4 I__236 (
            .O(N__1717),
            .I(\arse.seqcounterZ0Z_4 ));
    LocalMux I__235 (
            .O(N__1712),
            .I(\arse.seqcounterZ0Z_4 ));
    CascadeMux I__234 (
            .O(N__1707),
            .I(N__1703));
    InMux I__233 (
            .O(N__1706),
            .I(N__1700));
    InMux I__232 (
            .O(N__1703),
            .I(N__1697));
    LocalMux I__231 (
            .O(N__1700),
            .I(\arse.seqcounter_i_4 ));
    LocalMux I__230 (
            .O(N__1697),
            .I(\arse.seqcounter_i_4 ));
    InMux I__229 (
            .O(N__1692),
            .I(\arses.un2_counter_cry_1 ));
    InMux I__228 (
            .O(N__1689),
            .I(\arses.un2_counter_cry_2 ));
    InMux I__227 (
            .O(N__1686),
            .I(\arses.un2_counter_cry_3 ));
    InMux I__226 (
            .O(N__1683),
            .I(N__1679));
    InMux I__225 (
            .O(N__1682),
            .I(N__1676));
    LocalMux I__224 (
            .O(N__1679),
            .I(\arses.counterZ0Z_5 ));
    LocalMux I__223 (
            .O(N__1676),
            .I(\arses.counterZ0Z_5 ));
    InMux I__222 (
            .O(N__1671),
            .I(\arses.un2_counter_cry_4 ));
    InMux I__221 (
            .O(N__1668),
            .I(N__1664));
    InMux I__220 (
            .O(N__1667),
            .I(N__1661));
    LocalMux I__219 (
            .O(N__1664),
            .I(\arses.counterZ0Z_6 ));
    LocalMux I__218 (
            .O(N__1661),
            .I(\arses.counterZ0Z_6 ));
    InMux I__217 (
            .O(N__1656),
            .I(\arses.un2_counter_cry_5 ));
    InMux I__216 (
            .O(N__1653),
            .I(N__1649));
    InMux I__215 (
            .O(N__1652),
            .I(N__1646));
    LocalMux I__214 (
            .O(N__1649),
            .I(\arses.counterZ0Z_7 ));
    LocalMux I__213 (
            .O(N__1646),
            .I(\arses.counterZ0Z_7 ));
    InMux I__212 (
            .O(N__1641),
            .I(\arses.un2_counter_cry_6 ));
    CascadeMux I__211 (
            .O(N__1638),
            .I(\arse.divseven.N_65_i_cascade_ ));
    CascadeMux I__210 (
            .O(N__1635),
            .I(N__1626));
    InMux I__209 (
            .O(N__1634),
            .I(N__1623));
    InMux I__208 (
            .O(N__1633),
            .I(N__1620));
    InMux I__207 (
            .O(N__1632),
            .I(N__1617));
    InMux I__206 (
            .O(N__1631),
            .I(N__1614));
    InMux I__205 (
            .O(N__1630),
            .I(N__1607));
    InMux I__204 (
            .O(N__1629),
            .I(N__1607));
    InMux I__203 (
            .O(N__1626),
            .I(N__1607));
    LocalMux I__202 (
            .O(N__1623),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__201 (
            .O(N__1620),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__200 (
            .O(N__1617),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__199 (
            .O(N__1614),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__198 (
            .O(N__1607),
            .I(\arse.divseven.counterZ0Z_2 ));
    IoInMux I__197 (
            .O(N__1596),
            .I(N__1593));
    LocalMux I__196 (
            .O(N__1593),
            .I(N__1590));
    Odrv12 I__195 (
            .O(N__1590),
            .I(\arse.divseven.doutZ0Z_0 ));
    CEMux I__194 (
            .O(N__1587),
            .I(N__1583));
    CEMux I__193 (
            .O(N__1586),
            .I(N__1580));
    LocalMux I__192 (
            .O(N__1583),
            .I(N__1577));
    LocalMux I__191 (
            .O(N__1580),
            .I(N__1574));
    Span4Mux_h I__190 (
            .O(N__1577),
            .I(N__1569));
    Span4Mux_s3_v I__189 (
            .O(N__1574),
            .I(N__1569));
    Odrv4 I__188 (
            .O(N__1569),
            .I(\arse.divseven.N_65_i_0 ));
    InMux I__187 (
            .O(N__1566),
            .I(N__1563));
    LocalMux I__186 (
            .O(N__1563),
            .I(\arse.seqcounterZ0Z_0 ));
    InMux I__185 (
            .O(N__1560),
            .I(N__1557));
    LocalMux I__184 (
            .O(N__1557),
            .I(\arse.seqcounterZ0Z_1 ));
    InMux I__183 (
            .O(N__1554),
            .I(\arse.un1_seqcounter_1_cry_0 ));
    InMux I__182 (
            .O(N__1551),
            .I(N__1548));
    LocalMux I__181 (
            .O(N__1548),
            .I(\arse.seqcounterZ0Z_2 ));
    InMux I__180 (
            .O(N__1545),
            .I(\arse.un1_seqcounter_1_cry_1 ));
    InMux I__179 (
            .O(N__1542),
            .I(N__1539));
    LocalMux I__178 (
            .O(N__1539),
            .I(\arse.seqcounterZ1Z_3 ));
    InMux I__177 (
            .O(N__1536),
            .I(\arse.un1_seqcounter_1_cry_2 ));
    InMux I__176 (
            .O(N__1533),
            .I(\arse.un1_seqcounter_1_cry_3 ));
    CascadeMux I__175 (
            .O(N__1530),
            .I(\arse.divseven.N_60_i_cascade_ ));
    CEMux I__174 (
            .O(N__1527),
            .I(N__1524));
    LocalMux I__173 (
            .O(N__1524),
            .I(N__1521));
    Odrv12 I__172 (
            .O(N__1521),
            .I(\arse.divseven.counter_6_sqmuxa ));
    CascadeMux I__171 (
            .O(N__1518),
            .I(\arse.divseven.N_6_cascade_ ));
    CascadeMux I__170 (
            .O(N__1515),
            .I(\arse.divseven.un1_dout_2_sqmuxa_i_o2_0_cascade_ ));
    CascadeMux I__169 (
            .O(N__1512),
            .I(\arse.divseven.N_10_cascade_ ));
    InMux I__168 (
            .O(N__1509),
            .I(N__1504));
    InMux I__167 (
            .O(N__1508),
            .I(N__1501));
    InMux I__166 (
            .O(N__1507),
            .I(N__1495));
    LocalMux I__165 (
            .O(N__1504),
            .I(N__1490));
    LocalMux I__164 (
            .O(N__1501),
            .I(N__1490));
    InMux I__163 (
            .O(N__1500),
            .I(N__1487));
    InMux I__162 (
            .O(N__1499),
            .I(N__1482));
    InMux I__161 (
            .O(N__1498),
            .I(N__1482));
    LocalMux I__160 (
            .O(N__1495),
            .I(\arse.divseven.counterZ0Z_1 ));
    Odrv4 I__159 (
            .O(N__1490),
            .I(\arse.divseven.counterZ0Z_1 ));
    LocalMux I__158 (
            .O(N__1487),
            .I(\arse.divseven.counterZ0Z_1 ));
    LocalMux I__157 (
            .O(N__1482),
            .I(\arse.divseven.counterZ0Z_1 ));
    InMux I__156 (
            .O(N__1473),
            .I(N__1465));
    InMux I__155 (
            .O(N__1472),
            .I(N__1462));
    InMux I__154 (
            .O(N__1471),
            .I(N__1459));
    InMux I__153 (
            .O(N__1470),
            .I(N__1452));
    InMux I__152 (
            .O(N__1469),
            .I(N__1452));
    InMux I__151 (
            .O(N__1468),
            .I(N__1452));
    LocalMux I__150 (
            .O(N__1465),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__149 (
            .O(N__1462),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__148 (
            .O(N__1459),
            .I(\arse.divseven.counterZ0Z_0 ));
    LocalMux I__147 (
            .O(N__1452),
            .I(\arse.divseven.counterZ0Z_0 ));
    CascadeMux I__146 (
            .O(N__1443),
            .I(N__1439));
    CascadeMux I__145 (
            .O(N__1442),
            .I(N__1436));
    InMux I__144 (
            .O(N__1439),
            .I(N__1432));
    InMux I__143 (
            .O(N__1436),
            .I(N__1429));
    CascadeMux I__142 (
            .O(N__1435),
            .I(N__1426));
    LocalMux I__141 (
            .O(N__1432),
            .I(N__1418));
    LocalMux I__140 (
            .O(N__1429),
            .I(N__1418));
    InMux I__139 (
            .O(N__1426),
            .I(N__1415));
    InMux I__138 (
            .O(N__1425),
            .I(N__1412));
    InMux I__137 (
            .O(N__1424),
            .I(N__1407));
    InMux I__136 (
            .O(N__1423),
            .I(N__1407));
    Odrv4 I__135 (
            .O(N__1418),
            .I(\arse.divseven.sevenZ0 ));
    LocalMux I__134 (
            .O(N__1415),
            .I(\arse.divseven.sevenZ0 ));
    LocalMux I__133 (
            .O(N__1412),
            .I(\arse.divseven.sevenZ0 ));
    LocalMux I__132 (
            .O(N__1407),
            .I(\arse.divseven.sevenZ0 ));
    IoInMux I__131 (
            .O(N__1398),
            .I(N__1395));
    LocalMux I__130 (
            .O(N__1395),
            .I(N__1392));
    Odrv12 I__129 (
            .O(N__1392),
            .I(\arse.divseven.doutZ0Z_1 ));
    IoInMux I__128 (
            .O(N__1389),
            .I(N__1386));
    LocalMux I__127 (
            .O(N__1386),
            .I(N__1383));
    IoSpan4Mux I__126 (
            .O(N__1383),
            .I(N__1380));
    Span4Mux_s3_h I__125 (
            .O(N__1380),
            .I(N__1377));
    Sp12to4 I__124 (
            .O(N__1377),
            .I(N__1374));
    Span12Mux_v I__123 (
            .O(N__1374),
            .I(N__1371));
    Span12Mux_h I__122 (
            .O(N__1371),
            .I(N__1368));
    Odrv12 I__121 (
            .O(N__1368),
            .I(\top_pll_nrtthrth.PLLOUTCORE_0 ));
    INV \INVarse.diveight.dout_0C  (
            .O(\INVarse.diveight.dout_0C_net ),
            .I(N__2942));
    INV \INVarse.divseven.dout_nesr_0C  (
            .O(\INVarse.divseven.dout_nesr_0C_net ),
            .I(N__2940));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(\arses.un2_counter_cry_8 ),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    ICE_GB \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5  (
            .USERSIGNALTOGLOBALBUFFER(N__1389),
            .GLOBALBUFFEROUTPUT(PLLOUTCORE_0_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \arse.divseven.dout_esr_1_LC_4_4_6 .C_ON=1'b0;
    defparam \arse.divseven.dout_esr_1_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_esr_1_LC_4_4_6 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \arse.divseven.dout_esr_1_LC_4_4_6  (
            .in0(N__1634),
            .in1(N__1508),
            .in2(N__1443),
            .in3(N__1473),
            .lcout(\arse.divseven.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2936),
            .ce(N__1587),
            .sr(N__2879));
    defparam \arse.divseven.seven_RNO_0_LC_4_5_5 .C_ON=1'b0;
    defparam \arse.divseven.seven_RNO_0_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.seven_RNO_0_LC_4_5_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \arse.divseven.seven_RNO_0_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__1425),
            .in2(_gnd_net_),
            .in3(N__1471),
            .lcout(),
            .ltout(\arse.divseven.N_60_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.seven_RNO_LC_4_5_6 .C_ON=1'b0;
    defparam \arse.divseven.seven_RNO_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.seven_RNO_LC_4_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \arse.divseven.seven_RNO_LC_4_5_6  (
            .in0(N__1632),
            .in1(N__1500),
            .in2(N__1530),
            .in3(N__3130),
            .lcout(\arse.divseven.counter_6_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.seven_LC_4_6_0 .C_ON=1'b0;
    defparam \arse.divseven.seven_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.seven_LC_4_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \arse.divseven.seven_LC_4_6_0  (
            .in0(N__3372),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\arse.divseven.sevenZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2935),
            .ce(N__1527),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_ns_2_0__m5_LC_5_4_1 .C_ON=1'b0;
    defparam \arse.divseven.counter_ns_2_0__m5_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.counter_ns_2_0__m5_LC_5_4_1 .LUT_INIT=16'b0100110010110011;
    LogicCell40 \arse.divseven.counter_ns_2_0__m5_LC_5_4_1  (
            .in0(N__1633),
            .in1(N__1509),
            .in2(N__1442),
            .in3(N__1472),
            .lcout(),
            .ltout(\arse.divseven.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_1_LC_5_4_2 .C_ON=1'b0;
    defparam \arse.divseven.counter_1_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_1_LC_5_4_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \arse.divseven.counter_1_LC_5_4_2  (
            .in0(N__3125),
            .in1(_gnd_net_),
            .in2(N__1518),
            .in3(_gnd_net_),
            .lcout(\arse.divseven.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2939),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_ns_2_0__m3_s_LC_5_5_1 .C_ON=1'b0;
    defparam \arse.divseven.counter_ns_2_0__m3_s_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.counter_ns_2_0__m3_s_LC_5_5_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \arse.divseven.counter_ns_2_0__m3_s_LC_5_5_1  (
            .in0(N__1499),
            .in1(N__1424),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\arse.divseven.un1_dout_2_sqmuxa_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_0_LC_5_5_2 .C_ON=1'b0;
    defparam \arse.divseven.counter_0_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_0_LC_5_5_2 .LUT_INIT=16'b1001010100000000;
    LogicCell40 \arse.divseven.counter_0_LC_5_5_2  (
            .in0(N__1470),
            .in1(N__1630),
            .in2(N__1515),
            .in3(N__3097),
            .lcout(\arse.divseven.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2937),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_ns_2_0__m9_LC_5_5_3 .C_ON=1'b0;
    defparam \arse.divseven.counter_ns_2_0__m9_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.counter_ns_2_0__m9_LC_5_5_3 .LUT_INIT=16'b0001100111010101;
    LogicCell40 \arse.divseven.counter_ns_2_0__m9_LC_5_5_3  (
            .in0(N__1629),
            .in1(N__1507),
            .in2(N__1435),
            .in3(N__1469),
            .lcout(),
            .ltout(\arse.divseven.N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_2_LC_5_5_4 .C_ON=1'b0;
    defparam \arse.divseven.counter_2_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_2_LC_5_5_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \arse.divseven.counter_2_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1512),
            .in3(N__3096),
            .lcout(\arse.divseven.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2937),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_RNI8ECT_0_LC_5_5_5 .C_ON=1'b0;
    defparam \arse.divseven.counter_RNI8ECT_0_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.counter_RNI8ECT_0_LC_5_5_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \arse.divseven.counter_RNI8ECT_0_LC_5_5_5  (
            .in0(N__1498),
            .in1(N__1468),
            .in2(N__1635),
            .in3(N__1423),
            .lcout(),
            .ltout(\arse.divseven.N_65_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_RNI04101_0_LC_5_5_6 .C_ON=1'b0;
    defparam \arse.divseven.counter_RNI04101_0_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.counter_RNI04101_0_LC_5_5_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \arse.divseven.counter_RNI04101_0_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1638),
            .in3(N__2841),
            .lcout(\arse.divseven.N_65_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_nesr_0_LC_6_4_3 .C_ON=1'b0;
    defparam \arse.divseven.dout_nesr_0_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_nesr_0_LC_6_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.divseven.dout_nesr_0_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1631),
            .lcout(\arse.divseven.doutZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.divseven.dout_nesr_0C_net ),
            .ce(N__1586),
            .sr(N__2842));
    defparam \arse.seqreset_e_0_RNIOLK2_LC_6_5_5 .C_ON=1'b0;
    defparam \arse.seqreset_e_0_RNIOLK2_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \arse.seqreset_e_0_RNIOLK2_LC_6_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.seqreset_e_0_RNIOLK2_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3074),
            .lcout(\arse.seqreset_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqreset_e_0_LC_6_6_7 .C_ON=1'b0;
    defparam \arse.seqreset_e_0_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \arse.seqreset_e_0_LC_6_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.seqreset_e_0_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1725),
            .lcout(\arse.seqresetZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2938),
            .ce(N__2325),
            .sr(_gnd_net_));
    defparam \arse.seqcounter_0_LC_6_9_0 .C_ON=1'b1;
    defparam \arse.seqcounter_0_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \arse.seqcounter_0_LC_6_9_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \arse.seqcounter_0_LC_6_9_0  (
            .in0(N__2307),
            .in1(N__1566),
            .in2(N__1707),
            .in3(N__1706),
            .lcout(\arse.seqcounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\arse.un1_seqcounter_1_cry_0 ),
            .clk(N__2934),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqcounter_1_LC_6_9_1 .C_ON=1'b1;
    defparam \arse.seqcounter_1_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \arse.seqcounter_1_LC_6_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \arse.seqcounter_1_LC_6_9_1  (
            .in0(N__2309),
            .in1(N__1560),
            .in2(_gnd_net_),
            .in3(N__1554),
            .lcout(\arse.seqcounterZ0Z_1 ),
            .ltout(),
            .carryin(\arse.un1_seqcounter_1_cry_0 ),
            .carryout(\arse.un1_seqcounter_1_cry_1 ),
            .clk(N__2934),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqcounter_2_LC_6_9_2 .C_ON=1'b1;
    defparam \arse.seqcounter_2_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \arse.seqcounter_2_LC_6_9_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \arse.seqcounter_2_LC_6_9_2  (
            .in0(N__2308),
            .in1(N__1551),
            .in2(_gnd_net_),
            .in3(N__1545),
            .lcout(\arse.seqcounterZ0Z_2 ),
            .ltout(),
            .carryin(\arse.un1_seqcounter_1_cry_1 ),
            .carryout(\arse.un1_seqcounter_1_cry_2 ),
            .clk(N__2934),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqcounter_3_LC_6_9_3 .C_ON=1'b1;
    defparam \arse.seqcounter_3_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \arse.seqcounter_3_LC_6_9_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \arse.seqcounter_3_LC_6_9_3  (
            .in0(N__2310),
            .in1(N__1542),
            .in2(_gnd_net_),
            .in3(N__1536),
            .lcout(\arse.seqcounterZ1Z_3 ),
            .ltout(),
            .carryin(\arse.un1_seqcounter_1_cry_2 ),
            .carryout(\arse.un1_seqcounter_1_cry_3 ),
            .clk(N__2934),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqcounter_4_LC_6_9_4 .C_ON=1'b0;
    defparam \arse.seqcounter_4_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \arse.seqcounter_4_LC_6_9_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \arse.seqcounter_4_LC_6_9_4  (
            .in0(N__1721),
            .in1(N__2311),
            .in2(_gnd_net_),
            .in3(N__1533),
            .lcout(\arse.seqcounterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2934),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqcounter_RNIEP0A_4_LC_6_9_5 .C_ON=1'b0;
    defparam \arse.seqcounter_RNIEP0A_4_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \arse.seqcounter_RNIEP0A_4_LC_6_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.seqcounter_RNIEP0A_4_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1720),
            .lcout(\arse.seqcounter_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIA58_5_LC_9_3_0 .C_ON=1'b0;
    defparam \arses.counter_RNIA58_5_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIA58_5_LC_9_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \arses.counter_RNIA58_5_LC_9_3_0  (
            .in0(N__1652),
            .in1(N__1667),
            .in2(N__1782),
            .in3(N__1682),
            .lcout(\arses.un1_counterlto8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.un2_counter_cry_1_c_LC_9_4_0 .C_ON=1'b1;
    defparam \arses.un2_counter_cry_1_c_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \arses.un2_counter_cry_1_c_LC_9_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \arses.un2_counter_cry_1_c_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__1896),
            .in2(N__1875),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\arses.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_2_LC_9_4_1 .C_ON=1'b1;
    defparam \arses.counter_2_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_2_LC_9_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_2_LC_9_4_1  (
            .in0(N__2201),
            .in1(N__1932),
            .in2(_gnd_net_),
            .in3(N__1692),
            .lcout(\arses.counterZ0Z_2 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_1 ),
            .carryout(\arses.un2_counter_cry_2 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_3_LC_9_4_2 .C_ON=1'b1;
    defparam \arses.counter_3_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_3_LC_9_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_3_LC_9_4_2  (
            .in0(N__2193),
            .in1(N__1944),
            .in2(_gnd_net_),
            .in3(N__1689),
            .lcout(\arses.counterZ0Z_3 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_2 ),
            .carryout(\arses.un2_counter_cry_3 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_4_LC_9_4_3 .C_ON=1'b1;
    defparam \arses.counter_4_LC_9_4_3 .SEQ_MODE=4'b1001;
    defparam \arses.counter_4_LC_9_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_4_LC_9_4_3  (
            .in0(N__2202),
            .in1(N__1919),
            .in2(_gnd_net_),
            .in3(N__1686),
            .lcout(\arses.counterZ0Z_4 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_3 ),
            .carryout(\arses.un2_counter_cry_4 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_5_LC_9_4_4 .C_ON=1'b1;
    defparam \arses.counter_5_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_5_LC_9_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_5_LC_9_4_4  (
            .in0(N__2194),
            .in1(N__1683),
            .in2(_gnd_net_),
            .in3(N__1671),
            .lcout(\arses.counterZ0Z_5 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_4 ),
            .carryout(\arses.un2_counter_cry_5 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_6_LC_9_4_5 .C_ON=1'b1;
    defparam \arses.counter_6_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_6_LC_9_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_6_LC_9_4_5  (
            .in0(N__2203),
            .in1(N__1668),
            .in2(_gnd_net_),
            .in3(N__1656),
            .lcout(\arses.counterZ0Z_6 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_5 ),
            .carryout(\arses.un2_counter_cry_6 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_7_LC_9_4_6 .C_ON=1'b1;
    defparam \arses.counter_7_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \arses.counter_7_LC_9_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_7_LC_9_4_6  (
            .in0(N__2195),
            .in1(N__1653),
            .in2(_gnd_net_),
            .in3(N__1641),
            .lcout(\arses.counterZ0Z_7 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_6 ),
            .carryout(\arses.un2_counter_cry_7 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_8_LC_9_4_7 .C_ON=1'b1;
    defparam \arses.counter_8_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \arses.counter_8_LC_9_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_8_LC_9_4_7  (
            .in0(N__2204),
            .in1(N__1781),
            .in2(_gnd_net_),
            .in3(N__1767),
            .lcout(\arses.counterZ0Z_8 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_7 ),
            .carryout(\arses.un2_counter_cry_8 ),
            .clk(N__2473),
            .ce(),
            .sr(N__1852));
    defparam \arses.counter_9_LC_9_5_0 .C_ON=1'b1;
    defparam \arses.counter_9_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \arses.counter_9_LC_9_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_9_LC_9_5_0  (
            .in0(N__2192),
            .in1(N__1794),
            .in2(_gnd_net_),
            .in3(N__1764),
            .lcout(\arses.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\arses.un2_counter_cry_9 ),
            .clk(N__2474),
            .ce(),
            .sr(N__1854));
    defparam \arses.counter_10_LC_9_5_1 .C_ON=1'b1;
    defparam \arses.counter_10_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_10_LC_9_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_10_LC_9_5_1  (
            .in0(N__2198),
            .in1(N__1827),
            .in2(_gnd_net_),
            .in3(N__1761),
            .lcout(\arses.counterZ0Z_10 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_9 ),
            .carryout(\arses.un2_counter_cry_10 ),
            .clk(N__2474),
            .ce(),
            .sr(N__1854));
    defparam \arses.counter_11_LC_9_5_2 .C_ON=1'b1;
    defparam \arses.counter_11_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_11_LC_9_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_11_LC_9_5_2  (
            .in0(N__2190),
            .in1(N__1808),
            .in2(_gnd_net_),
            .in3(N__1758),
            .lcout(\arses.counterZ0Z_11 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_10 ),
            .carryout(\arses.un2_counter_cry_11 ),
            .clk(N__2474),
            .ce(),
            .sr(N__1854));
    defparam \arses.counter_12_LC_9_5_3 .C_ON=1'b1;
    defparam \arses.counter_12_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \arses.counter_12_LC_9_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_12_LC_9_5_3  (
            .in0(N__2199),
            .in1(N__2040),
            .in2(_gnd_net_),
            .in3(N__1755),
            .lcout(\arses.counterZ0Z_12 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_11 ),
            .carryout(\arses.un2_counter_cry_12 ),
            .clk(N__2474),
            .ce(),
            .sr(N__1854));
    defparam \arses.counter_13_LC_9_5_4 .C_ON=1'b1;
    defparam \arses.counter_13_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_13_LC_9_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_13_LC_9_5_4  (
            .in0(N__2191),
            .in1(N__2055),
            .in2(_gnd_net_),
            .in3(N__1752),
            .lcout(\arses.counterZ0Z_13 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_12 ),
            .carryout(\arses.un2_counter_cry_13 ),
            .clk(N__2474),
            .ce(),
            .sr(N__1854));
    defparam \arses.counter_14_LC_9_5_5 .C_ON=1'b0;
    defparam \arses.counter_14_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_14_LC_9_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_14_LC_9_5_5  (
            .in0(N__2200),
            .in1(N__2067),
            .in2(_gnd_net_),
            .in3(N__1749),
            .lcout(\arses.counterZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2474),
            .ce(),
            .sr(N__1854));
    defparam masterreset_ibuf_RNIKP26_LC_9_6_2.C_ON=1'b0;
    defparam masterreset_ibuf_RNIKP26_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam masterreset_ibuf_RNIKP26_LC_9_6_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 masterreset_ibuf_RNIKP26_LC_9_6_2 (
            .in0(N__2326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(masterreset_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_0_LC_10_1_0 .C_ON=1'b0;
    defparam \arse.diveight.dout_0_LC_10_1_0 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_0_LC_10_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.diveight.dout_0_LC_10_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2981),
            .lcout(\arse.diveight.doutZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.diveight.dout_0C_net ),
            .ce(),
            .sr(N__2887));
    defparam \arse.diveight.counter_2_LC_10_3_3 .C_ON=1'b0;
    defparam \arse.diveight.counter_2_LC_10_3_3 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_2_LC_10_3_3 .LUT_INIT=16'b0110110000000000;
    LogicCell40 \arse.diveight.counter_2_LC_10_3_3  (
            .in0(N__1961),
            .in1(N__2977),
            .in2(N__1974),
            .in3(N__3139),
            .lcout(\arse.diveight.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2941),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_1_LC_10_3_6 .C_ON=1'b0;
    defparam \arse.diveight.counter_1_LC_10_3_6 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_1_LC_10_3_6 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \arse.diveight.counter_1_LC_10_3_6  (
            .in0(_gnd_net_),
            .in1(N__3137),
            .in2(N__1962),
            .in3(N__1970),
            .lcout(\arse.diveight.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2941),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_0_LC_10_3_7 .C_ON=1'b0;
    defparam \arse.diveight.counter_0_LC_10_3_7 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_0_LC_10_3_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \arse.diveight.counter_0_LC_10_3_7  (
            .in0(N__3138),
            .in1(N__1957),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\arse.diveight.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2941),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI1L5_2_LC_10_4_0 .C_ON=1'b0;
    defparam \arses.counter_RNI1L5_2_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI1L5_2_LC_10_4_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \arses.counter_RNI1L5_2_LC_10_4_0  (
            .in0(N__1943),
            .in1(N__1931),
            .in2(_gnd_net_),
            .in3(N__1890),
            .lcout(),
            .ltout(\arses.un1_counterlto4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOKH_1_LC_10_4_1 .C_ON=1'b0;
    defparam \arses.counter_RNIOKH_1_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOKH_1_LC_10_4_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \arses.counter_RNIOKH_1_LC_10_4_1  (
            .in0(N__1920),
            .in1(N__1867),
            .in2(N__1905),
            .in3(N__1902),
            .lcout(\arses.un1_counterlt11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_0_LC_10_4_3 .C_ON=1'b0;
    defparam \arses.counter_0_LC_10_4_3 .SEQ_MODE=4'b1001;
    defparam \arses.counter_0_LC_10_4_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \arses.counter_0_LC_10_4_3  (
            .in0(N__1891),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2197),
            .lcout(\arses.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2471),
            .ce(),
            .sr(N__1853));
    defparam \arses.counter_1_LC_10_4_4 .C_ON=1'b0;
    defparam \arses.counter_1_LC_10_4_4 .SEQ_MODE=4'b1001;
    defparam \arses.counter_1_LC_10_4_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \arses.counter_1_LC_10_4_4  (
            .in0(N__2196),
            .in1(_gnd_net_),
            .in2(N__1874),
            .in3(N__1892),
            .lcout(\arses.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2471),
            .ce(),
            .sr(N__1853));
    defparam \arses.counter_RNI04C4_9_LC_10_5_2 .C_ON=1'b0;
    defparam \arses.counter_RNI04C4_9_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI04C4_9_LC_10_5_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \arses.counter_RNI04C4_9_LC_10_5_2  (
            .in0(N__1826),
            .in1(N__1815),
            .in2(N__1809),
            .in3(N__1793),
            .lcout(),
            .ltout(\arses.un1_counterlt13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOS0A_14_LC_10_5_3 .C_ON=1'b0;
    defparam \arses.counter_RNIOS0A_14_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOS0A_14_LC_10_5_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \arses.counter_RNIOS0A_14_LC_10_5_3  (
            .in0(N__2066),
            .in1(N__2054),
            .in2(N__2043),
            .in3(N__2039),
            .lcout(\arses.counter8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_4_LC_11_3_0 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_4_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_4_LC_11_3_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \debounceconsolereset.counter_4_LC_11_3_0  (
            .in0(N__2552),
            .in1(N__2358),
            .in2(N__2598),
            .in3(N__2375),
            .lcout(\debounceconsolereset.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2469),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_2_LC_11_3_2 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_2_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_2_LC_11_3_2 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \debounceconsolereset.counter_2_LC_11_3_2  (
            .in0(N__2550),
            .in1(N__2007),
            .in2(N__2028),
            .in3(N__2596),
            .lcout(\debounceconsolereset.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2469),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_RNO_1_LC_11_3_4 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNO_1_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNO_1_LC_11_3_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \debounceconsolereset.out_RNO_1_LC_11_3_4  (
            .in0(N__2024),
            .in1(N__2374),
            .in2(N__1997),
            .in3(N__2520),
            .lcout(\debounceconsolereset.out_cnv_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNISLFD_2_LC_11_3_5 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_RNISLFD_2_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNISLFD_2_LC_11_3_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \debounceconsolereset.counter_RNISLFD_2_LC_11_3_5  (
            .in0(N__2373),
            .in1(N__1989),
            .in2(_gnd_net_),
            .in3(N__2023),
            .lcout(\debounceconsolereset.un1_counterlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_3_LC_11_3_6 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_3_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_3_LC_11_3_6 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \debounceconsolereset.counter_3_LC_11_3_6  (
            .in0(N__2551),
            .in1(N__2385),
            .in2(N__1998),
            .in3(N__2597),
            .lcout(\debounceconsolereset.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2469),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_0_LC_11_3_7 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_0_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_0_LC_11_3_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \debounceconsolereset.counter_0_LC_11_3_7  (
            .in0(N__2521),
            .in1(N__2591),
            .in2(_gnd_net_),
            .in3(N__2553),
            .lcout(\debounceconsolereset.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2469),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_11_4_0 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_1_c_LC_11_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_1_c_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__2491),
            .in2(N__2525),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\debounceconsolereset.un3_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_11_4_1 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_11_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__2022),
            .in2(_gnd_net_),
            .in3(N__2001),
            .lcout(\debounceconsolereset.un3_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_1 ),
            .carryout(\debounceconsolereset.un3_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_11_4_2 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_11_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(N__1996),
            .in2(_gnd_net_),
            .in3(N__2379),
            .lcout(\debounceconsolereset.un3_counter_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_2 ),
            .carryout(\debounceconsolereset.un3_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_3_THRU_LUT4_0_LC_11_4_3 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_3_THRU_LUT4_0_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_3_THRU_LUT4_0_LC_11_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_3_THRU_LUT4_0_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__2376),
            .in2(_gnd_net_),
            .in3(N__2352),
            .lcout(\debounceconsolereset.un3_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_3 ),
            .carryout(\debounceconsolereset.un3_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_cry_4_THRU_LUT4_0_LC_11_4_4 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_cry_4_THRU_LUT4_0_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_cry_4_THRU_LUT4_0_LC_11_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounceconsolereset.un3_counter_cry_4_THRU_LUT4_0_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__2110),
            .in2(_gnd_net_),
            .in3(N__2349),
            .lcout(\debounceconsolereset.un3_counter_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_cry_4 ),
            .carryout(\debounceconsolereset.un3_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_6_LC_11_4_5 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_6_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_6_LC_11_4_5 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \debounceconsolereset.counter_6_LC_11_4_5  (
            .in0(N__2085),
            .in1(N__2595),
            .in2(N__2559),
            .in3(N__2346),
            .lcout(\debounceconsolereset.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2470),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_LC_11_4_6 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_LC_11_4_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \arses.clock_out_RNIR6ER_LC_11_4_6  (
            .in0(N__2334),
            .in1(N__2132),
            .in2(_gnd_net_),
            .in3(N__2189),
            .lcout(clock_out_RNIR6ER),
            .ltout(clock_out_RNIR6ER_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNI4RTH1_6_LC_11_4_7 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_RNI4RTH1_6_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNI4RTH1_6_LC_11_4_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \debounceconsolereset.counter_RNI4RTH1_6_LC_11_4_7  (
            .in0(N__2109),
            .in1(N__2083),
            .in2(N__2343),
            .in3(N__2340),
            .lcout(\debounceconsolereset.counter_RNI4RTH1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_LC_11_5_1 .C_ON=1'b0;
    defparam \arses.clock_out_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \arses.clock_out_LC_11_5_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \arses.clock_out_LC_11_5_1  (
            .in0(N__2333),
            .in1(N__2133),
            .in2(_gnd_net_),
            .in3(N__2205),
            .lcout(\arses.clock_out_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2472),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_5_LC_11_5_2 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_5_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_5_LC_11_5_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \debounceconsolereset.counter_5_LC_11_5_2  (
            .in0(N__2554),
            .in1(N__2112),
            .in2(N__2121),
            .in3(N__2590),
            .lcout(\debounceconsolereset.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2472),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_RNO_0_LC_11_5_5 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNO_0_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNO_0_LC_11_5_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \debounceconsolereset.out_RNO_0_LC_11_5_5  (
            .in0(N__2111),
            .in1(N__2094),
            .in2(N__2498),
            .in3(N__2084),
            .lcout(),
            .ltout(\debounceconsolereset.out_cnv_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_LC_11_5_6 .C_ON=1'b0;
    defparam \debounceconsolereset.out_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.out_LC_11_5_6 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \debounceconsolereset.out_LC_11_5_6  (
            .in0(N__2616),
            .in1(N__2589),
            .in2(N__2601),
            .in3(N__3239),
            .lcout(apureset_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2472),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_1_LC_11_5_7 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_1_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_1_LC_11_5_7 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \debounceconsolereset.counter_1_LC_11_5_7  (
            .in0(N__2588),
            .in1(N__2555),
            .in2(N__2499),
            .in3(N__2526),
            .lcout(\debounceconsolereset.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2472),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.counter_1_LC_15_5_3 .C_ON=1'b0;
    defparam \arse.arse.counter_1_LC_15_5_3 .SEQ_MODE=4'b1001;
    defparam \arse.arse.counter_1_LC_15_5_3 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \arse.arse.counter_1_LC_15_5_3  (
            .in0(N__2726),
            .in1(N__2433),
            .in2(N__2409),
            .in3(N__2670),
            .lcout(\arse.arse.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2943),
            .ce(),
            .sr(N__2866));
    defparam \arse.arse.counter_2_LC_15_5_7 .C_ON=1'b0;
    defparam \arse.arse.counter_2_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \arse.arse.counter_2_LC_15_5_7 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \arse.arse.counter_2_LC_15_5_7  (
            .in0(N__2727),
            .in1(N__2810),
            .in2(N__2787),
            .in3(N__2671),
            .lcout(\arse.arse.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2943),
            .ce(),
            .sr(N__2866));
    defparam \arse.arse.counter_RNIHKTF1_1_LC_15_6_3 .C_ON=1'b0;
    defparam \arse.arse.counter_RNIHKTF1_1_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \arse.arse.counter_RNIHKTF1_1_LC_15_6_3 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \arse.arse.counter_RNIHKTF1_1_LC_15_6_3  (
            .in0(N__2808),
            .in1(N__2401),
            .in2(_gnd_net_),
            .in3(N__2430),
            .lcout(\arse.un1_counterlt4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_5.C_ON=1'b0;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2478),
            .lcout(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.counter_0_LC_16_5_4 .C_ON=1'b0;
    defparam \arse.arse.counter_0_LC_16_5_4 .SEQ_MODE=4'b1001;
    defparam \arse.arse.counter_0_LC_16_5_4 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \arse.arse.counter_0_LC_16_5_4  (
            .in0(N__2811),
            .in1(N__2716),
            .in2(_gnd_net_),
            .in3(N__2432),
            .lcout(\arse.arse.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2945),
            .ce(),
            .sr(N__2880));
    defparam \arse.arse.counter_3_LC_16_5_6 .C_ON=1'b0;
    defparam \arse.arse.counter_3_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \arse.arse.counter_3_LC_16_5_6 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \arse.arse.counter_3_LC_16_5_6  (
            .in0(N__2717),
            .in1(N__2748),
            .in2(N__2775),
            .in3(N__2675),
            .lcout(\arse.arse.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2945),
            .ce(),
            .sr(N__2880));
    defparam \arse.arse.un16_counter_cry_1_c_LC_16_6_0 .C_ON=1'b1;
    defparam \arse.arse.un16_counter_cry_1_c_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \arse.arse.un16_counter_cry_1_c_LC_16_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \arse.arse.un16_counter_cry_1_c_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__2431),
            .in2(N__2408),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\arse.arse.un16_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.un16_counter_cry_1_THRU_LUT4_0_LC_16_6_1 .C_ON=1'b1;
    defparam \arse.arse.un16_counter_cry_1_THRU_LUT4_0_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \arse.arse.un16_counter_cry_1_THRU_LUT4_0_LC_16_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.arse.un16_counter_cry_1_THRU_LUT4_0_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(N__2809),
            .in2(_gnd_net_),
            .in3(N__2778),
            .lcout(\arse.arse.un16_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\arse.arse.un16_counter_cry_1 ),
            .carryout(\arse.arse.un16_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.un16_counter_cry_2_THRU_LUT4_0_LC_16_6_2 .C_ON=1'b1;
    defparam \arse.arse.un16_counter_cry_2_THRU_LUT4_0_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \arse.arse.un16_counter_cry_2_THRU_LUT4_0_LC_16_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.arse.un16_counter_cry_2_THRU_LUT4_0_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__2747),
            .in2(_gnd_net_),
            .in3(N__2766),
            .lcout(\arse.arse.un16_counter_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\arse.arse.un16_counter_cry_2 ),
            .carryout(\arse.arse.un16_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.counter_4_LC_16_6_3 .C_ON=1'b0;
    defparam \arse.arse.counter_4_LC_16_6_3 .SEQ_MODE=4'b1001;
    defparam \arse.arse.counter_4_LC_16_6_3 .LUT_INIT=16'b0101000110100010;
    LogicCell40 \arse.arse.counter_4_LC_16_6_3  (
            .in0(N__2760),
            .in1(N__2715),
            .in2(N__2682),
            .in3(N__2763),
            .lcout(\arse.arse.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2944),
            .ce(),
            .sr(N__2888));
    defparam \arse.arse.counter_RNIRIUV_4_LC_17_6_0 .C_ON=1'b0;
    defparam \arse.arse.counter_RNIRIUV_4_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \arse.arse.counter_RNIRIUV_4_LC_17_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.arse.counter_RNIRIUV_4_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__2759),
            .in2(_gnd_net_),
            .in3(N__2746),
            .lcout(\arse.un1_counterlto4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.ddd.Q_esr_RNO_LC_18_5_2 .C_ON=1'b0;
    defparam \arse.ddd.Q_esr_RNO_LC_18_5_2 .SEQ_MODE=4'b0000;
    defparam \arse.ddd.Q_esr_RNO_LC_18_5_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \arse.ddd.Q_esr_RNO_LC_18_5_2  (
            .in0(_gnd_net_),
            .in1(N__3284),
            .in2(_gnd_net_),
            .in3(N__2622),
            .lcout(\arse.ddd.N_33_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.clock_out_RNIM09F_LC_18_6_2 .C_ON=1'b0;
    defparam \arse.arse.clock_out_RNIM09F_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \arse.arse.clock_out_RNIM09F_LC_18_6_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \arse.arse.clock_out_RNIM09F_LC_18_6_2  (
            .in0(_gnd_net_),
            .in1(N__3269),
            .in2(_gnd_net_),
            .in3(N__2632),
            .lcout(),
            .ltout(\arse.G_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.seqreset_e_0_RNIQTP13_LC_18_6_3 .C_ON=1'b0;
    defparam \arse.seqreset_e_0_RNIQTP13_LC_18_6_3 .SEQ_MODE=4'b0000;
    defparam \arse.seqreset_e_0_RNIQTP13_LC_18_6_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \arse.seqreset_e_0_RNIQTP13_LC_18_6_3  (
            .in0(N__2713),
            .in1(N__2677),
            .in2(N__2730),
            .in3(N__3127),
            .lcout(\arse.seqreset_e_0_RNIQTPZ0Z13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.arse.clock_out_LC_18_6_5 .C_ON=1'b0;
    defparam \arse.arse.clock_out_LC_18_6_5 .SEQ_MODE=4'b1000;
    defparam \arse.arse.clock_out_LC_18_6_5 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \arse.arse.clock_out_LC_18_6_5  (
            .in0(N__2714),
            .in1(N__2678),
            .in2(N__2640),
            .in3(N__3128),
            .lcout(\arse.clock_out_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2946),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.ddd.Q_esr_RNO_0_LC_18_6_7 .C_ON=1'b0;
    defparam \arse.ddd.Q_esr_RNO_0_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \arse.ddd.Q_esr_RNO_0_LC_18_6_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \arse.ddd.Q_esr_RNO_0_LC_18_6_7  (
            .in0(N__2712),
            .in1(N__2676),
            .in2(N__2639),
            .in3(N__3126),
            .lcout(\arse.ddd.Q_esr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_18_16_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_16_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_16_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.ddd.Q_esr_LC_19_5_1 .C_ON=1'b0;
    defparam \arse.ddd.Q_esr_LC_19_5_1 .SEQ_MODE=4'b1000;
    defparam \arse.ddd.Q_esr_LC_19_5_1 .LUT_INIT=16'b1000000010100000;
    LogicCell40 \arse.ddd.Q_esr_LC_19_5_1  (
            .in0(N__3255),
            .in1(N__3218),
            .in2(N__3146),
            .in3(N__3206),
            .lcout(cpureset_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2947),
            .ce(N__3297),
            .sr(N__3291));
    defparam \arse.l2.un1_Q_LC_19_6_1 .C_ON=1'b0;
    defparam \arse.l2.un1_Q_LC_19_6_1 .SEQ_MODE=4'b0000;
    defparam \arse.l2.un1_Q_LC_19_6_1 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \arse.l2.un1_Q_LC_19_6_1  (
            .in0(N__3219),
            .in1(N__3207),
            .in2(N__3273),
            .in3(N__3129),
            .lcout(G_73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.l1.N_23_0_i_LC_20_4_4 .C_ON=1'b0;
    defparam \arse.l1.N_23_0_i_LC_20_4_4 .SEQ_MODE=4'b0000;
    defparam \arse.l1.N_23_0_i_LC_20_4_4 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \arse.l1.N_23_0_i_LC_20_4_4  (
            .in0(N__3036),
            .in1(N__3199),
            .in2(N__3164),
            .in3(N__3147),
            .lcout(G_74),
            .ltout(G_74_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.io_0_RNIIG08_LC_20_4_5 .C_ON=1'b0;
    defparam \arse.divseven.io_0_RNIIG08_LC_20_4_5 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.io_0_RNIIG08_LC_20_4_5 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \arse.divseven.io_0_RNIIG08_LC_20_4_5  (
            .in0(N__3030),
            .in1(_gnd_net_),
            .in2(N__3018),
            .in3(_gnd_net_),
            .lcout(arse_un1_apuclk_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_1_LC_30_5_5 .C_ON=1'b0;
    defparam \arse.diveight.dout_1_LC_30_5_5 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_1_LC_30_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.diveight.dout_1_LC_30_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2994),
            .lcout(\arse.diveight.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2948),
            .ce(),
            .sr(N__2892));
endmodule // top
