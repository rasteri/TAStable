-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 12 2024 12:32:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    masterreset : in std_logic;
    led4 : out std_logic;
    lcol3 : out std_logic;
    led5 : out std_logic;
    lcol2 : out std_logic;
    led6 : out std_logic;
    led2 : out std_logic;
    lcol1 : out std_logic;
    deldn : in std_logic;
    cpuclk : out std_logic;
    apureset : out std_logic;
    altreset : in std_logic;
    led7 : out std_logic;
    led3 : out std_logic;
    lcol4 : out std_logic;
    delup : in std_logic;
    cpureset : out std_logic;
    apusync : in std_logic;
    PACKAGEPIN : in std_logic;
    led8 : out std_logic;
    led1 : out std_logic;
    consolereset : in std_logic;
    apuclk : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \arse.un1_io_0_1_g\ : std_logic;
signal \top_pll_nrtthrth.PLLOUTCORE\ : std_logic;
signal \arse.divseven.io_0_D_IN_0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal masterreset_c_i : std_logic;
signal \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\ : std_logic;
signal deldn_c : std_logic;
signal leds_1_i_1 : std_logic;
signal leds_1_i_3 : std_logic;
signal \dig2.leds_cnst_2_cascade_\ : std_logic;
signal leds_1_i_2 : std_logic;
signal \olddnZ0\ : std_logic;
signal debounceddn : std_logic;
signal \dig2.un1_leds114_0\ : std_logic;
signal \dig2.i2_mux_cascade_\ : std_logic;
signal \dig2.leds_cnst_1\ : std_logic;
signal \dig2.m29_bm_0_cascade_\ : std_logic;
signal \dig2.m30_ns_1\ : std_logic;
signal \dig2.m23_am_0\ : std_logic;
signal \dig2.m29_am_0\ : std_logic;
signal \dig2.N_38\ : std_logic;
signal \dig2.m23_bm_0\ : std_logic;
signal \dig2.m34_am_0_cascade_\ : std_logic;
signal \dig2.m34_bm_0\ : std_logic;
signal \dig2.N_35\ : std_logic;
signal \delayConstant16_i_cascade_\ : std_logic;
signal \oldupZ0\ : std_logic;
signal \un1_delayConstant_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_21_11_0_\ : std_logic;
signal \olddn_RNISQ7L1Z0Z_2\ : std_logic;
signal \un1_delayConstant_cry_0\ : std_logic;
signal \olddn_RNISQ7L1Z0Z_0\ : std_logic;
signal \un1_delayConstant_cry_1\ : std_logic;
signal \olddn_RNISQ7L1Z0Z_3\ : std_logic;
signal \un1_delayConstant_cry_2\ : std_logic;
signal \olddn_RNISQ7L1Z0Z_1\ : std_logic;
signal \un1_delayConstant_cry_3\ : std_logic;
signal \olddn_RNISQ7LZ0Z1\ : std_logic;
signal \un1_delayConstant_cry_4\ : std_logic;
signal \olddn_RNISQ7L1Z0Z_4\ : std_logic;
signal \un1_delayConstant_cry_5\ : std_logic;
signal \un1_delayConstant_cry_6\ : std_logic;
signal \delayConstant16_i\ : std_logic;
signal \olddn_RNI1J1RZ0\ : std_logic;
signal \delayConstantZ0Z_6\ : std_logic;
signal \dig2.m8_am_0_cascade_\ : std_logic;
signal \dig2.N_9\ : std_logic;
signal \slowclk_0_cascade_\ : std_logic;
signal slowclk_0 : std_logic;
signal \delayConstantZ0Z_4\ : std_logic;
signal \delayConstantZ0Z_5\ : std_logic;
signal \dig2.m8_bm_0\ : std_logic;
signal col_1_1 : std_logic;
signal \col_1_1_cascade_\ : std_logic;
signal \dig1.m34_am_cascade_\ : std_logic;
signal \dig1.m34_bm\ : std_logic;
signal \bfn_22_8_0_\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_1\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_2\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_3\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_2_THRU_CO\ : std_logic;
signal \debounceconsolereset.un3_counter_cry_1_THRU_CO\ : std_logic;
signal \clock_out_RNIR6ER_0_cascade_\ : std_logic;
signal \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_\ : std_logic;
signal \debounceconsolereset.counter_RNINST81Z0Z_4\ : std_logic;
signal masterreset_c : std_logic;
signal slowclk : std_logic;
signal debouncedn_counter_4 : std_logic;
signal debouncedn_counter_1 : std_logic;
signal debouncedn_counter_0 : std_logic;
signal debouncedn_counter_2 : std_logic;
signal \debouncedn.out_cnvZ0Z_1\ : std_logic;
signal debouncedn_counter_3 : std_logic;
signal consolereset_c : std_logic;
signal altreset_c : std_logic;
signal \out_cnv_cascade_\ : std_logic;
signal \un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2\ : std_logic;
signal \un1_delayConstant_cry_3_0_c_RNITFZ0Z062\ : std_logic;
signal \un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2\ : std_logic;
signal \un1_delayConstant_cry_1_0_c_RNIP5KDZ0Z2\ : std_logic;
signal \dig1.m8_am_cascade_\ : std_logic;
signal \dig1.m8_bm\ : std_logic;
signal \dig1.N_9_cascade_\ : std_logic;
signal \dig1.i2_mux\ : std_logic;
signal \dig1.m23_bm\ : std_logic;
signal \dig1.m29_bm_cascade_\ : std_logic;
signal \dig1.m23_am\ : std_logic;
signal \dig1.m29_am_cascade_\ : std_logic;
signal \dig1.m30_ns_1\ : std_logic;
signal \delayConstantZ0Z_0\ : std_logic;
signal \delayConstantZ0Z_2\ : std_logic;
signal \dig1.leds_cnst_1\ : std_logic;
signal leds_1_i_0_1 : std_logic;
signal \dig1.N_38\ : std_logic;
signal \dig1.N_35\ : std_logic;
signal leds_1_i_0_3 : std_logic;
signal \dig1.un1_leds114_0\ : std_logic;
signal \dig1.leds_cnst_2\ : std_logic;
signal leds_1_i_0_2 : std_logic;
signal lcol1_c : std_logic;
signal lcol2_c : std_logic;
signal lcol3_c : std_logic;
signal \colZ0Z_1\ : std_logic;
signal \colZ0Z_0\ : std_logic;
signal lcol4_c : std_logic;
signal \clock_out_RNIR6ER_0\ : std_logic;
signal \INVarse.doingsevenC_net\ : std_logic;
signal \delayConstant_fastZ0Z_2\ : std_logic;
signal \delayConstant_fastZ0Z_0\ : std_logic;
signal \arse.g0_3_cascade_\ : std_logic;
signal \arse.g0_7_cascade_\ : std_logic;
signal \arse.cpuresetoutreg_1_sqmuxa_cascade_\ : std_logic;
signal \arse.cpuresetoutregZ0\ : std_logic;
signal \INVarse.cpuresetoutregC_net\ : std_logic;
signal \arses.un1_counterlto8_2_cascade_\ : std_logic;
signal \arses.un1_counterlto4_2\ : std_logic;
signal \arses.un1_counterlt11_cascade_\ : std_logic;
signal \arses.un1_counterlt13_0_cascade_\ : std_logic;
signal \arses.counterZ0Z_0\ : std_logic;
signal \arses.counterZ0Z_1\ : std_logic;
signal \bfn_23_10_0_\ : std_logic;
signal \arses.counterZ0Z_2\ : std_logic;
signal \arses.un2_counter_cry_1\ : std_logic;
signal \arses.counterZ0Z_3\ : std_logic;
signal \arses.un2_counter_cry_2\ : std_logic;
signal \arses.counterZ0Z_4\ : std_logic;
signal \arses.un2_counter_cry_3\ : std_logic;
signal \arses.counterZ0Z_5\ : std_logic;
signal \arses.un2_counter_cry_4\ : std_logic;
signal \arses.counterZ0Z_6\ : std_logic;
signal \arses.un2_counter_cry_5\ : std_logic;
signal \arses.counterZ0Z_7\ : std_logic;
signal \arses.un2_counter_cry_6\ : std_logic;
signal \arses.counterZ0Z_8\ : std_logic;
signal \arses.un2_counter_cry_7\ : std_logic;
signal \arses.un2_counter_cry_8\ : std_logic;
signal \arses.counterZ0Z_9\ : std_logic;
signal \bfn_23_11_0_\ : std_logic;
signal \arses.counterZ0Z_10\ : std_logic;
signal \arses.un2_counter_cry_9\ : std_logic;
signal \arses.counterZ0Z_11\ : std_logic;
signal \arses.un2_counter_cry_10\ : std_logic;
signal \arses.counterZ0Z_12\ : std_logic;
signal \arses.un2_counter_cry_11\ : std_logic;
signal \arses.counterZ0Z_13\ : std_logic;
signal \arses.un2_counter_cry_12\ : std_logic;
signal \arses.counter8\ : std_logic;
signal \arses.un2_counter_cry_13\ : std_logic;
signal \arses.counterZ0Z_14\ : std_logic;
signal masterreset_c_i_g : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \arse.doingseven3\ : std_logic;
signal \arse.g0_i_a3_4_cascade_\ : std_logic;
signal \arse.N_6\ : std_logic;
signal \arse.doingseven3_6\ : std_logic;
signal \arse.doingseven3_1\ : std_logic;
signal \arse.doingseven3_6_cascade_\ : std_logic;
signal \arse.cpuresetcountZ0Z_0\ : std_logic;
signal \bfn_24_8_0_\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_0\ : std_logic;
signal \arse.cpuresetcountZ0Z_2\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_1\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_2\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_3\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_4\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_5\ : std_logic;
signal \arse.un1_cpuresetcount_1_cry_6\ : std_logic;
signal \INVarse.cpuresetcount_0C_net\ : std_logic;
signal \delayConstantZ0Z_7\ : std_logic;
signal \arse.cpuresetcountZ0Z_1\ : std_logic;
signal \delayConstantZ0Z_1\ : std_logic;
signal \arse.cpuresetcountZ0Z_7\ : std_logic;
signal \arse.g0_1\ : std_logic;
signal \delayConstant_fastZ0Z_6\ : std_logic;
signal \delayConstant_fastZ0Z_5\ : std_logic;
signal \arse.cpuresetcountZ0Z_6\ : std_logic;
signal \arse.cpuresetcountZ0Z_5\ : std_logic;
signal \arse.g0_4\ : std_logic;
signal \delayConstant_fastZ0Z_4\ : std_logic;
signal \delayConstantZ0Z_3\ : std_logic;
signal \arse.cpuresetcountZ0Z_4\ : std_logic;
signal \arse.cpuresetcountZ0Z_3\ : std_logic;
signal \arse.g0_2\ : std_logic;
signal \arse.doingsevenZ0\ : std_logic;
signal \arse.divseven.N_41_0\ : std_logic;
signal delup_c : std_logic;
signal debouncedup : std_logic;
signal \PACKAGEPIN_0_c_g\ : std_logic;
signal out_cnv : std_logic;
signal \arse.divseven.dout_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \arse.divseven.doutZ0Z_0\ : std_logic;
signal \INVarse.divseven.dout_0C_net\ : std_logic;
signal \arse.divseven.counterZ0Z_1\ : std_logic;
signal \arse.divseven.sevenZ0\ : std_logic;
signal \arse.doingseven4\ : std_logic;
signal \INVarse.cpuclkresetC_net\ : std_logic;
signal debouncedconsolereset_i : std_logic;
signal apusync_c : std_logic;
signal \arse.apusynclatchedZ0\ : std_logic;
signal \INVarse.apusynclatchedC_net\ : std_logic;
signal \arse.diveight.counterZ0Z_0\ : std_logic;
signal \arse.diveight.counterZ0Z_1\ : std_logic;
signal \arse.diveight.doutZ0Z_1\ : std_logic;
signal \arse.cpuclkresetZ0\ : std_logic;
signal \arse.diveight.counterZ0Z_2\ : std_logic;
signal \arse.diveight.doutZ1Z_0\ : std_logic;
signal debouncedconsolereset : std_logic;
signal \arse.apuresetoutregZ0\ : std_logic;
signal \INVarse.diveight.dout_0C_net\ : std_logic;
signal \arse.divseven.counterZ0Z_2\ : std_logic;
signal \arse.divseven.un1_dout_2_sqmuxa_0_o3_0\ : std_logic;
signal \arse.divseven.counterZ0Z_0\ : std_logic;
signal \arse.divseven.doutZ0Z_1\ : std_logic;
signal \PLLOUTCORE_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PACKAGEPIN_wire\ : std_logic;
signal masterreset_wire : std_logic;
signal led3_wire : std_logic;
signal apuclk_wire : std_logic;
signal cpureset_wire : std_logic;
signal lcol3_wire : std_logic;
signal deldn_wire : std_logic;
signal led2_wire : std_logic;
signal delup_wire : std_logic;
signal led6_wire : std_logic;
signal led8_wire : std_logic;
signal altreset_wire : std_logic;
signal led4_wire : std_logic;
signal apureset_wire : std_logic;
signal lcol4_wire : std_logic;
signal cpuclk_wire : std_logic;
signal led5_wire : std_logic;
signal consolereset_wire : std_logic;
signal lcol2_wire : std_logic;
signal led1_wire : std_logic;
signal apusync_wire : std_logic;
signal led7_wire : std_logic;
signal lcol1_wire : std_logic;
signal \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \PACKAGEPIN_wire\ <= PACKAGEPIN;
    masterreset_wire <= masterreset;
    led3 <= led3_wire;
    apuclk <= apuclk_wire;
    cpureset <= cpureset_wire;
    lcol3 <= lcol3_wire;
    deldn_wire <= deldn;
    led2 <= led2_wire;
    delup_wire <= delup;
    led6 <= led6_wire;
    led8 <= led8_wire;
    altreset_wire <= altreset;
    led4 <= led4_wire;
    apureset <= apureset_wire;
    lcol4 <= lcol4_wire;
    cpuclk <= cpuclk_wire;
    led5 <= led5_wire;
    consolereset_wire <= consolereset;
    lcol2 <= lcol2_wire;
    led1 <= led1_wire;
    apusync_wire <= apusync;
    led7 <= led7_wire;
    lcol1 <= lcol1_wire;
    \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_nrtthrth.top_pll_nrtthrth_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "010",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \top_pll_nrtthrth.PLLOUTCORE\,
            REFERENCECLK => \N__2337\,
            RESETB => \N__3213\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \top_pll_nrtthrth.top_pll_nrtthrth_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PACKAGEPIN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5959\,
            GLOBALBUFFEROUTPUT => \PACKAGEPIN_0_c_g\
        );

    \PACKAGEPIN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5961\,
            DIN => \N__5960\,
            DOUT => \N__5959\,
            PACKAGEPIN => \PACKAGEPIN_wire\
        );

    \PACKAGEPIN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5961\,
            PADOUT => \N__5960\,
            PADIN => \N__5959\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \masterreset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5950\,
            DIN => \N__5949\,
            DOUT => \N__5948\,
            PACKAGEPIN => masterreset_wire
        );

    \masterreset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5950\,
            PADOUT => \N__5949\,
            PADIN => \N__5948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => masterreset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5941\,
            DIN => \N__5940\,
            DOUT => \N__5939\,
            PACKAGEPIN => led3_wire
        );

    \led3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5941\,
            PADOUT => \N__5940\,
            PADIN => \N__5939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.divseven.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5932\,
            DIN => \N__5931\,
            DOUT => \N__5930\,
            PACKAGEPIN => apuclk_wire
        );

    \arse.divseven.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5932\,
            PADOUT => \N__5931\,
            PADIN => \N__5930\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__5411\,
            OUTPUTENABLE => \N__4415\,
            DIN0 => \arse.divseven.io_0_D_IN_0\,
            DOUT0 => \N__5217\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5395\
        );

    \arse.io_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5923\,
            DIN => \N__5922\,
            DOUT => \N__5921\,
            PACKAGEPIN => cpureset_wire
        );

    \arse.io_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5923\,
            PADOUT => \N__5922\,
            PADIN => \N__5921\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4206\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5400\
        );

    \lcol3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5914\,
            DIN => \N__5913\,
            DOUT => \N__5912\,
            PACKAGEPIN => lcol3_wire
        );

    \lcol3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5914\,
            PADOUT => \N__5913\,
            PADIN => \N__5912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3978\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \deldn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5905\,
            DIN => \N__5904\,
            DOUT => \N__5903\,
            PACKAGEPIN => deldn_wire
        );

    \deldn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5905\,
            PADOUT => \N__5904\,
            PADIN => \N__5903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => deldn_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5896\,
            DIN => \N__5895\,
            DOUT => \N__5894\,
            PACKAGEPIN => led2_wire
        );

    \led2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5896\,
            PADOUT => \N__5895\,
            PADIN => \N__5894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3324\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delup_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5887\,
            DIN => \N__5886\,
            DOUT => \N__5885\,
            PACKAGEPIN => delup_wire
        );

    \delup_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5887\,
            PADOUT => \N__5886\,
            PADIN => \N__5885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delup_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led6_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5878\,
            DIN => \N__5877\,
            DOUT => \N__5876\,
            PACKAGEPIN => led6_wire
        );

    \led6_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5878\,
            PADOUT => \N__5877\,
            PADIN => \N__5876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led8_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5869\,
            DIN => \N__5868\,
            DOUT => \N__5867\,
            PACKAGEPIN => led8_wire
        );

    \led8_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5869\,
            PADOUT => \N__5868\,
            PADIN => \N__5867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \altreset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5860\,
            DIN => \N__5859\,
            DOUT => \N__5858\,
            PACKAGEPIN => altreset_wire
        );

    \altreset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5860\,
            PADOUT => \N__5859\,
            PADIN => \N__5858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => altreset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5851\,
            DIN => \N__5850\,
            DOUT => \N__5849\,
            PACKAGEPIN => led4_wire
        );

    \led4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5851\,
            PADOUT => \N__5850\,
            PADIN => \N__5849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4086\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5842\,
            DIN => \N__5841\,
            DOUT => \N__5840\,
            PACKAGEPIN => apureset_wire
        );

    \arse.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "010101",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5842\,
            PADOUT => \N__5841\,
            PADIN => \N__5840\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5508\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5399\
        );

    \lcol4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5833\,
            DIN => \N__5832\,
            DOUT => \N__5831\,
            PACKAGEPIN => lcol4_wire
        );

    \lcol4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5833\,
            PADOUT => \N__5832\,
            PADIN => \N__5831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \arse.diveight.io_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5824\,
            DIN => \N__5823\,
            DOUT => \N__5822\,
            PACKAGEPIN => cpuclk_wire
        );

    \arse.diveight.io_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "100001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5824\,
            PADOUT => \N__5823\,
            PADIN => \N__5822\,
            CLOCKENABLE => 'H',
            DOUT1 => \N__5628\,
            OUTPUTENABLE => \N__4422\,
            DIN0 => OPEN,
            DOUT0 => \N__5562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => \N__5399\
        );

    \led5_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5815\,
            DIN => \N__5814\,
            DOUT => \N__5813\,
            PACKAGEPIN => led5_wire
        );

    \led5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5815\,
            PADOUT => \N__5814\,
            PADIN => \N__5813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \consolereset_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5806\,
            DIN => \N__5805\,
            DOUT => \N__5804\,
            PACKAGEPIN => consolereset_wire
        );

    \consolereset_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5806\,
            PADOUT => \N__5805\,
            PADIN => \N__5804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => consolereset_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5797\,
            DIN => \N__5796\,
            DOUT => \N__5795\,
            PACKAGEPIN => lcol2_wire
        );

    \lcol2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5797\,
            PADOUT => \N__5796\,
            PADIN => \N__5795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5788\,
            DIN => \N__5787\,
            DOUT => \N__5786\,
            PACKAGEPIN => led1_wire
        );

    \led1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5788\,
            PADOUT => \N__5787\,
            PADIN => \N__5786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4393\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \apusync_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5779\,
            DIN => \N__5778\,
            DOUT => \N__5777\,
            PACKAGEPIN => apusync_wire
        );

    \apusync_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5779\,
            PADOUT => \N__5778\,
            PADIN => \N__5777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => apusync_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5770\,
            DIN => \N__5769\,
            DOUT => \N__5768\,
            PACKAGEPIN => led7_wire
        );

    \led7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5770\,
            PADOUT => \N__5769\,
            PADIN => \N__5768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2442\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \lcol1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5761\,
            DIN => \N__5760\,
            DOUT => \N__5759\,
            PACKAGEPIN => lcol1_wire
        );

    \lcol1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5761\,
            PADOUT => \N__5760\,
            PADIN => \N__5759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1368\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5739\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5736\
        );

    \I__1366\ : Span12Mux_v
    port map (
            O => \N__5736\,
            I => \N__5733\
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__5733\,
            I => apusync_c
        );

    \I__1364\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5726\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__5729\,
            I => \N__5721\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__5726\,
            I => \N__5718\
        );

    \I__1361\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5715\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5712\
        );

    \I__1359\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5709\
        );

    \I__1358\ : Span4Mux_v
    port map (
            O => \N__5718\,
            I => \N__5704\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5704\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__5712\,
            I => \N__5699\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__5709\,
            I => \N__5699\
        );

    \I__1354\ : Span4Mux_v
    port map (
            O => \N__5704\,
            I => \N__5693\
        );

    \I__1353\ : Span4Mux_v
    port map (
            O => \N__5699\,
            I => \N__5693\
        );

    \I__1352\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5690\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__5693\,
            I => \N__5685\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__5690\,
            I => \N__5685\
        );

    \I__1349\ : Span4Mux_h
    port map (
            O => \N__5685\,
            I => \N__5681\
        );

    \I__1348\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5678\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__5681\,
            I => \arse.apusynclatchedZ0\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__5678\,
            I => \arse.apusynclatchedZ0\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__5673\,
            I => \N__5668\
        );

    \I__1344\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5664\
        );

    \I__1343\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5661\
        );

    \I__1342\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5656\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5656\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5664\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5661\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__5656\,
            I => \arse.diveight.counterZ0Z_0\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__5649\,
            I => \N__5645\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__5648\,
            I => \N__5642\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5638\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5633\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5633\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__5638\,
            I => \arse.diveight.counterZ0Z_1\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__5633\,
            I => \arse.diveight.counterZ0Z_1\
        );

    \I__1330\ : IoInMux
    port map (
            O => \N__5628\,
            I => \N__5625\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__5625\,
            I => \arse.diveight.doutZ0Z_1\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5618\
        );

    \I__1327\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5615\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5611\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__5615\,
            I => \N__5608\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5602\
        );

    \I__1323\ : Span4Mux_s1_h
    port map (
            O => \N__5611\,
            I => \N__5599\
        );

    \I__1322\ : Span4Mux_s1_h
    port map (
            O => \N__5608\,
            I => \N__5596\
        );

    \I__1321\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5589\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5589\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5589\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5602\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1317\ : Odrv4
    port map (
            O => \N__5599\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__5596\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__5589\,
            I => \arse.cpuclkresetZ0\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5575\
        );

    \I__1313\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5572\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5569\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5575\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__5572\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5569\,
            I => \arse.diveight.counterZ0Z_2\
        );

    \I__1308\ : IoInMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5559\,
            I => \arse.diveight.doutZ1Z_0\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5552\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5549\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5545\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5549\,
            I => \N__5542\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5539\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__5545\,
            I => \N__5536\
        );

    \I__1300\ : Span4Mux_s3_h
    port map (
            O => \N__5542\,
            I => \N__5531\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5539\,
            I => \N__5531\
        );

    \I__1298\ : Sp12to4
    port map (
            O => \N__5536\,
            I => \N__5528\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__5531\,
            I => \N__5525\
        );

    \I__1296\ : Span12Mux_s10_h
    port map (
            O => \N__5528\,
            I => \N__5521\
        );

    \I__1295\ : Sp12to4
    port map (
            O => \N__5525\,
            I => \N__5518\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5515\
        );

    \I__1293\ : Odrv12
    port map (
            O => \N__5521\,
            I => debouncedconsolereset
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__5518\,
            I => debouncedconsolereset
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5515\,
            I => debouncedconsolereset
        );

    \I__1290\ : IoInMux
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5505\,
            I => \arse.apuresetoutregZ0\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5499\,
            I => \N__5496\
        );

    \I__1286\ : Span4Mux_s1_h
    port map (
            O => \N__5496\,
            I => \N__5493\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__5493\,
            I => \N__5484\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5475\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5475\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5475\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5475\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5470\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5470\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__5484\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5475\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5470\,
            I => \arse.divseven.counterZ0Z_2\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__5463\,
            I => \N__5460\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5457\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5457\,
            I => \N__5454\
        );

    \I__1272\ : Span4Mux_s0_h
    port map (
            O => \N__5454\,
            I => \N__5451\
        );

    \I__1271\ : Span4Mux_h
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__5448\,
            I => \arse.divseven.un1_dout_2_sqmuxa_0_o3_0\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__1267\ : Span12Mux_v
    port map (
            O => \N__5439\,
            I => \N__5431\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5422\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5422\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5422\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5422\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5419\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__5431\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5422\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5419\,
            I => \arse.divseven.counterZ0Z_0\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5408\
        );

    \I__1257\ : IoInMux
    port map (
            O => \N__5411\,
            I => \N__5405\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5408\,
            I => \arse.divseven.doutZ0Z_1\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5405\,
            I => \arse.divseven.doutZ0Z_1\
        );

    \I__1254\ : ClkMux
    port map (
            O => \N__5400\,
            I => \N__5358\
        );

    \I__1253\ : ClkMux
    port map (
            O => \N__5399\,
            I => \N__5358\
        );

    \I__1252\ : ClkMux
    port map (
            O => \N__5398\,
            I => \N__5358\
        );

    \I__1251\ : ClkMux
    port map (
            O => \N__5397\,
            I => \N__5358\
        );

    \I__1250\ : ClkMux
    port map (
            O => \N__5396\,
            I => \N__5358\
        );

    \I__1249\ : ClkMux
    port map (
            O => \N__5395\,
            I => \N__5358\
        );

    \I__1248\ : ClkMux
    port map (
            O => \N__5394\,
            I => \N__5358\
        );

    \I__1247\ : ClkMux
    port map (
            O => \N__5393\,
            I => \N__5358\
        );

    \I__1246\ : ClkMux
    port map (
            O => \N__5392\,
            I => \N__5358\
        );

    \I__1245\ : ClkMux
    port map (
            O => \N__5391\,
            I => \N__5358\
        );

    \I__1244\ : ClkMux
    port map (
            O => \N__5390\,
            I => \N__5358\
        );

    \I__1243\ : ClkMux
    port map (
            O => \N__5389\,
            I => \N__5358\
        );

    \I__1242\ : ClkMux
    port map (
            O => \N__5388\,
            I => \N__5358\
        );

    \I__1241\ : ClkMux
    port map (
            O => \N__5387\,
            I => \N__5358\
        );

    \I__1240\ : GlobalMux
    port map (
            O => \N__5358\,
            I => \N__5355\
        );

    \I__1239\ : gio2CtrlBuf
    port map (
            O => \N__5355\,
            I => \PLLOUTCORE_g\
        );

    \I__1238\ : CEMux
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5346\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__5346\,
            I => \N__5343\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__5343\,
            I => \arse.divseven.N_41_0\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__1232\ : Span12Mux_v
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__1231\ : Odrv12
    port map (
            O => \N__5331\,
            I => delup_c
        );

    \I__1230\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5322\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5322\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5319\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__5319\,
            I => debouncedup
        );

    \I__1226\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5313\,
            I => \N__5290\
        );

    \I__1224\ : ClkMux
    port map (
            O => \N__5312\,
            I => \N__5247\
        );

    \I__1223\ : ClkMux
    port map (
            O => \N__5311\,
            I => \N__5247\
        );

    \I__1222\ : ClkMux
    port map (
            O => \N__5310\,
            I => \N__5247\
        );

    \I__1221\ : ClkMux
    port map (
            O => \N__5309\,
            I => \N__5247\
        );

    \I__1220\ : ClkMux
    port map (
            O => \N__5308\,
            I => \N__5247\
        );

    \I__1219\ : ClkMux
    port map (
            O => \N__5307\,
            I => \N__5247\
        );

    \I__1218\ : ClkMux
    port map (
            O => \N__5306\,
            I => \N__5247\
        );

    \I__1217\ : ClkMux
    port map (
            O => \N__5305\,
            I => \N__5247\
        );

    \I__1216\ : ClkMux
    port map (
            O => \N__5304\,
            I => \N__5247\
        );

    \I__1215\ : ClkMux
    port map (
            O => \N__5303\,
            I => \N__5247\
        );

    \I__1214\ : ClkMux
    port map (
            O => \N__5302\,
            I => \N__5247\
        );

    \I__1213\ : ClkMux
    port map (
            O => \N__5301\,
            I => \N__5247\
        );

    \I__1212\ : ClkMux
    port map (
            O => \N__5300\,
            I => \N__5247\
        );

    \I__1211\ : ClkMux
    port map (
            O => \N__5299\,
            I => \N__5247\
        );

    \I__1210\ : ClkMux
    port map (
            O => \N__5298\,
            I => \N__5247\
        );

    \I__1209\ : ClkMux
    port map (
            O => \N__5297\,
            I => \N__5247\
        );

    \I__1208\ : ClkMux
    port map (
            O => \N__5296\,
            I => \N__5247\
        );

    \I__1207\ : ClkMux
    port map (
            O => \N__5295\,
            I => \N__5247\
        );

    \I__1206\ : ClkMux
    port map (
            O => \N__5294\,
            I => \N__5247\
        );

    \I__1205\ : ClkMux
    port map (
            O => \N__5293\,
            I => \N__5247\
        );

    \I__1204\ : Glb2LocalMux
    port map (
            O => \N__5290\,
            I => \N__5247\
        );

    \I__1203\ : GlobalMux
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__1202\ : gio2CtrlBuf
    port map (
            O => \N__5244\,
            I => \PACKAGEPIN_0_c_g\
        );

    \I__1201\ : CEMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5234\
        );

    \I__1199\ : CEMux
    port map (
            O => \N__5237\,
            I => \N__5231\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__5234\,
            I => \N__5228\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5225\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__5228\,
            I => out_cnv
        );

    \I__1195\ : Odrv12
    port map (
            O => \N__5225\,
            I => out_cnv
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__5220\,
            I => \arse.divseven.dout_RNO_0Z0Z_0_cascade_\
        );

    \I__1193\ : IoInMux
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__1191\ : IoSpan4Mux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__1190\ : Span4Mux_s1_h
    port map (
            O => \N__5208\,
            I => \N__5204\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5201\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__5204\,
            I => \arse.divseven.doutZ0Z_0\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5201\,
            I => \arse.divseven.doutZ0Z_0\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__5196\,
            I => \N__5191\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__5195\,
            I => \N__5188\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__5194\,
            I => \N__5182\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5173\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5173\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5173\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5173\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5168\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5168\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5173\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5168\,
            I => \arse.divseven.counterZ0Z_1\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__5163\,
            I => \N__5158\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__5162\,
            I => \N__5154\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5143\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5143\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5143\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5143\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5138\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5138\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5143\,
            I => \arse.divseven.sevenZ0\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5138\,
            I => \arse.divseven.sevenZ0\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5127\
        );

    \I__1163\ : Odrv12
    port map (
            O => \N__5127\,
            I => \arse.doingseven4\
        );

    \I__1162\ : SRMux
    port map (
            O => \N__5124\,
            I => \N__5119\
        );

    \I__1161\ : SRMux
    port map (
            O => \N__5123\,
            I => \N__5116\
        );

    \I__1160\ : SRMux
    port map (
            O => \N__5122\,
            I => \N__5112\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5109\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5106\
        );

    \I__1157\ : SRMux
    port map (
            O => \N__5115\,
            I => \N__5103\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5112\,
            I => \N__5100\
        );

    \I__1155\ : Span4Mux_h
    port map (
            O => \N__5109\,
            I => \N__5097\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__5106\,
            I => \N__5092\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5103\,
            I => \N__5092\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__5100\,
            I => \N__5089\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__5097\,
            I => \N__5082\
        );

    \I__1150\ : Span4Mux_h
    port map (
            O => \N__5092\,
            I => \N__5082\
        );

    \I__1149\ : Span4Mux_v
    port map (
            O => \N__5089\,
            I => \N__5082\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__5082\,
            I => debouncedconsolereset_i
        );

    \I__1147\ : InMux
    port map (
            O => \N__5079\,
            I => \arse.un1_cpuresetcount_1_cry_6\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__5076\,
            I => \N__5072\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5067\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5064\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5071\,
            I => \N__5061\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__5070\,
            I => \N__5057\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5053\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5064\,
            I => \N__5050\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5061\,
            I => \N__5047\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5044\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5039\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5039\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__5053\,
            I => \N__5032\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__5050\,
            I => \N__5032\
        );

    \I__1133\ : Span4Mux_h
    port map (
            O => \N__5047\,
            I => \N__5032\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5044\,
            I => \delayConstantZ0Z_7\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5039\,
            I => \delayConstantZ0Z_7\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__5032\,
            I => \delayConstantZ0Z_7\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5019\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5016\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5013\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5008\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5008\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5016\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5013\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5008\,
            I => \arse.cpuresetcountZ0Z_1\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__1120\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4990\
        );

    \I__1119\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4983\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4983\
        );

    \I__1117\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4983\
        );

    \I__1116\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4974\
        );

    \I__1115\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4974\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__4990\,
            I => \N__4971\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__4983\,
            I => \N__4968\
        );

    \I__1112\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4961\
        );

    \I__1111\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4961\
        );

    \I__1110\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4961\
        );

    \I__1109\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4956\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4953\
        );

    \I__1107\ : Span4Mux_h
    port map (
            O => \N__4971\,
            I => \N__4946\
        );

    \I__1106\ : Span4Mux_v
    port map (
            O => \N__4968\,
            I => \N__4946\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__4961\,
            I => \N__4946\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4941\
        );

    \I__1103\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4941\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__4956\,
            I => \delayConstantZ0Z_1\
        );

    \I__1101\ : Odrv12
    port map (
            O => \N__4953\,
            I => \delayConstantZ0Z_1\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__4946\,
            I => \delayConstantZ0Z_1\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__4941\,
            I => \delayConstantZ0Z_1\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__4932\,
            I => \N__4926\
        );

    \I__1097\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4923\
        );

    \I__1096\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4920\
        );

    \I__1095\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4917\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4914\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__4923\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__4920\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4917\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__4914\,
            I => \arse.cpuresetcountZ0Z_7\
        );

    \I__1089\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4902\,
            I => \arse.g0_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__4893\,
            I => \N__4890\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__4890\,
            I => \delayConstant_fastZ0Z_6\
        );

    \I__1083\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__1081\ : Span4Mux_h
    port map (
            O => \N__4881\,
            I => \N__4878\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__4878\,
            I => \delayConstant_fastZ0Z_5\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__4875\,
            I => \N__4871\
        );

    \I__1078\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4866\
        );

    \I__1077\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4863\
        );

    \I__1076\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4858\
        );

    \I__1075\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4858\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__4866\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__4863\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4858\,
            I => \arse.cpuresetcountZ0Z_6\
        );

    \I__1071\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4845\
        );

    \I__1070\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4840\
        );

    \I__1069\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4840\
        );

    \I__1068\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4837\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__4845\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__4840\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__4837\,
            I => \arse.cpuresetcountZ0Z_5\
        );

    \I__1064\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__4827\,
            I => \arse.g0_4\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4821\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__4815\,
            I => \delayConstant_fastZ0Z_4\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__4812\,
            I => \N__4808\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4805\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4802\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4796\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4792\
        );

    \I__1053\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4789\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4784\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4784\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__4796\,
            I => \N__4781\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4778\
        );

    \I__1048\ : Span4Mux_v
    port map (
            O => \N__4792\,
            I => \N__4771\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4789\,
            I => \N__4771\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4784\,
            I => \N__4771\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__4781\,
            I => \delayConstantZ0Z_3\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4778\,
            I => \delayConstantZ0Z_3\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__4771\,
            I => \delayConstantZ0Z_3\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__4764\,
            I => \N__4760\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4755\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4752\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4747\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4747\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4755\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4752\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4747\,
            I => \arse.cpuresetcountZ0Z_4\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4733\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4726\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4726\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4726\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4723\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4733\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4726\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__4723\,
            I => \arse.cpuresetcountZ0Z_3\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4713\,
            I => \arse.g0_2\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4706\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4703\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4700\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4703\,
            I => \arse.doingsevenZ0\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__4700\,
            I => \arse.doingsevenZ0\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__4695\,
            I => \N__4692\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4689\,
            I => \arse.doingseven3_6\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4680\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4680\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4680\,
            I => \arse.doingseven3_1\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__4677\,
            I => \arse.doingseven3_6_cascade_\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4665\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4662\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4657\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4657\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4665\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4662\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4657\,
            I => \arse.cpuresetcountZ0Z_0\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4650\,
            I => \arse.un1_cpuresetcount_1_cry_0\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4639\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4639\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4636\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4633\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4639\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4636\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4633\,
            I => \arse.cpuresetcountZ0Z_2\
        );

    \I__996\ : InMux
    port map (
            O => \N__4626\,
            I => \arse.un1_cpuresetcount_1_cry_1\
        );

    \I__995\ : InMux
    port map (
            O => \N__4623\,
            I => \arse.un1_cpuresetcount_1_cry_2\
        );

    \I__994\ : InMux
    port map (
            O => \N__4620\,
            I => \arse.un1_cpuresetcount_1_cry_3\
        );

    \I__993\ : InMux
    port map (
            O => \N__4617\,
            I => \arse.un1_cpuresetcount_1_cry_4\
        );

    \I__992\ : InMux
    port map (
            O => \N__4614\,
            I => \arse.un1_cpuresetcount_1_cry_5\
        );

    \I__991\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4607\
        );

    \I__990\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4604\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4601\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4604\,
            I => \arses.counterZ0Z_11\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__4601\,
            I => \arses.counterZ0Z_11\
        );

    \I__986\ : InMux
    port map (
            O => \N__4596\,
            I => \arses.un2_counter_cry_10\
        );

    \I__985\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4589\
        );

    \I__984\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4586\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4589\,
            I => \N__4583\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4586\,
            I => \arses.counterZ0Z_12\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__4583\,
            I => \arses.counterZ0Z_12\
        );

    \I__980\ : InMux
    port map (
            O => \N__4578\,
            I => \arses.un2_counter_cry_11\
        );

    \I__979\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4571\
        );

    \I__978\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4568\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4571\,
            I => \N__4565\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4568\,
            I => \arses.counterZ0Z_13\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__4565\,
            I => \arses.counterZ0Z_13\
        );

    \I__974\ : InMux
    port map (
            O => \N__4560\,
            I => \arses.un2_counter_cry_12\
        );

    \I__973\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4542\
        );

    \I__972\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4539\
        );

    \I__971\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4536\
        );

    \I__970\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4524\
        );

    \I__969\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4524\
        );

    \I__968\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4524\
        );

    \I__967\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4524\
        );

    \I__966\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4517\
        );

    \I__965\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4517\
        );

    \I__964\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4517\
        );

    \I__963\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4510\
        );

    \I__962\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4510\
        );

    \I__961\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4510\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4542\,
            I => \N__4507\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4539\,
            I => \N__4502\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4502\
        );

    \I__957\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4493\
        );

    \I__956\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4493\
        );

    \I__955\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4493\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4486\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4486\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4510\,
            I => \N__4486\
        );

    \I__951\ : Span4Mux_h
    port map (
            O => \N__4507\,
            I => \N__4481\
        );

    \I__950\ : Span4Mux_v
    port map (
            O => \N__4502\,
            I => \N__4481\
        );

    \I__949\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4476\
        );

    \I__948\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4476\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4493\,
            I => \arses.counter8\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__4486\,
            I => \arses.counter8\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__4481\,
            I => \arses.counter8\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4476\,
            I => \arses.counter8\
        );

    \I__943\ : InMux
    port map (
            O => \N__4467\,
            I => \arses.un2_counter_cry_13\
        );

    \I__942\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4461\,
            I => \N__4457\
        );

    \I__940\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4454\
        );

    \I__939\ : Span4Mux_h
    port map (
            O => \N__4457\,
            I => \N__4451\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4454\,
            I => \arses.counterZ0Z_14\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__4451\,
            I => \arses.counterZ0Z_14\
        );

    \I__936\ : SRMux
    port map (
            O => \N__4446\,
            I => \N__4428\
        );

    \I__935\ : SRMux
    port map (
            O => \N__4445\,
            I => \N__4428\
        );

    \I__934\ : SRMux
    port map (
            O => \N__4444\,
            I => \N__4428\
        );

    \I__933\ : SRMux
    port map (
            O => \N__4443\,
            I => \N__4428\
        );

    \I__932\ : SRMux
    port map (
            O => \N__4442\,
            I => \N__4428\
        );

    \I__931\ : SRMux
    port map (
            O => \N__4441\,
            I => \N__4428\
        );

    \I__930\ : GlobalMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__929\ : gio2CtrlBuf
    port map (
            O => \N__4425\,
            I => masterreset_c_i_g
        );

    \I__928\ : IoInMux
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__926\ : IoSpan4Mux
    port map (
            O => \N__4416\,
            I => \N__4412\
        );

    \I__925\ : IoInMux
    port map (
            O => \N__4415\,
            I => \N__4409\
        );

    \I__924\ : IoSpan4Mux
    port map (
            O => \N__4412\,
            I => \N__4404\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4404\
        );

    \I__922\ : Span4Mux_s2_h
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__921\ : Span4Mux_h
    port map (
            O => \N__4401\,
            I => \N__4397\
        );

    \I__920\ : IoInMux
    port map (
            O => \N__4400\,
            I => \N__4394\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__4397\,
            I => \N__4390\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4394\,
            I => \N__4387\
        );

    \I__917\ : IoInMux
    port map (
            O => \N__4393\,
            I => \N__4384\
        );

    \I__916\ : Span12Mux_v
    port map (
            O => \N__4390\,
            I => \N__4381\
        );

    \I__915\ : Span4Mux_s1_v
    port map (
            O => \N__4387\,
            I => \N__4378\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4384\,
            I => \N__4375\
        );

    \I__913\ : Span12Mux_v
    port map (
            O => \N__4381\,
            I => \N__4372\
        );

    \I__912\ : Span4Mux_h
    port map (
            O => \N__4378\,
            I => \N__4369\
        );

    \I__911\ : Span12Mux_s1_v
    port map (
            O => \N__4375\,
            I => \N__4366\
        );

    \I__910\ : Odrv12
    port map (
            O => \N__4372\,
            I => \CONSTANT_ONE_NET\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4369\,
            I => \CONSTANT_ONE_NET\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__4366\,
            I => \CONSTANT_ONE_NET\
        );

    \I__907\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4356\,
            I => \arse.doingseven3\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4353\,
            I => \arse.g0_i_a3_4_cascade_\
        );

    \I__904\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4347\,
            I => \arse.N_6\
        );

    \I__902\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4340\
        );

    \I__901\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4337\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4340\,
            I => \arses.counterZ0Z_3\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4337\,
            I => \arses.counterZ0Z_3\
        );

    \I__898\ : InMux
    port map (
            O => \N__4332\,
            I => \arses.un2_counter_cry_2\
        );

    \I__897\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4325\
        );

    \I__896\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4322\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4325\,
            I => \arses.counterZ0Z_4\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4322\,
            I => \arses.counterZ0Z_4\
        );

    \I__893\ : InMux
    port map (
            O => \N__4317\,
            I => \arses.un2_counter_cry_3\
        );

    \I__892\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4310\
        );

    \I__891\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4307\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4310\,
            I => \arses.counterZ0Z_5\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4307\,
            I => \arses.counterZ0Z_5\
        );

    \I__888\ : InMux
    port map (
            O => \N__4302\,
            I => \arses.un2_counter_cry_4\
        );

    \I__887\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4295\
        );

    \I__886\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4292\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4295\,
            I => \arses.counterZ0Z_6\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4292\,
            I => \arses.counterZ0Z_6\
        );

    \I__883\ : InMux
    port map (
            O => \N__4287\,
            I => \arses.un2_counter_cry_5\
        );

    \I__882\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4280\
        );

    \I__881\ : InMux
    port map (
            O => \N__4283\,
            I => \N__4277\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4280\,
            I => \arses.counterZ0Z_7\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4277\,
            I => \arses.counterZ0Z_7\
        );

    \I__878\ : InMux
    port map (
            O => \N__4272\,
            I => \arses.un2_counter_cry_6\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4269\,
            I => \N__4265\
        );

    \I__876\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4262\
        );

    \I__875\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4259\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4262\,
            I => \arses.counterZ0Z_8\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4259\,
            I => \arses.counterZ0Z_8\
        );

    \I__872\ : InMux
    port map (
            O => \N__4254\,
            I => \arses.un2_counter_cry_7\
        );

    \I__871\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4247\
        );

    \I__870\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4244\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4247\,
            I => \N__4241\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4244\,
            I => \arses.counterZ0Z_9\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__4241\,
            I => \arses.counterZ0Z_9\
        );

    \I__866\ : InMux
    port map (
            O => \N__4236\,
            I => \bfn_23_11_0_\
        );

    \I__865\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4229\
        );

    \I__864\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4226\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4229\,
            I => \N__4223\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4226\,
            I => \arses.counterZ0Z_10\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__4223\,
            I => \arses.counterZ0Z_10\
        );

    \I__860\ : InMux
    port map (
            O => \N__4218\,
            I => \arses.un2_counter_cry_9\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \arse.g0_3_cascade_\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__4212\,
            I => \arse.g0_7_cascade_\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__4209\,
            I => \arse.cpuresetoutreg_1_sqmuxa_cascade_\
        );

    \I__856\ : IoInMux
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__854\ : Span4Mux_s0_h
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__853\ : Span4Mux_h
    port map (
            O => \N__4197\,
            I => \N__4193\
        );

    \I__852\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4190\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__4193\,
            I => \N__4187\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4190\,
            I => \arse.cpuresetoutregZ0\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__4187\,
            I => \arse.cpuresetoutregZ0\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__4182\,
            I => \arses.un1_counterlto8_2_cascade_\
        );

    \I__847\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4176\,
            I => \arses.un1_counterlto4_2\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4173\,
            I => \arses.un1_counterlt11_cascade_\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__4170\,
            I => \arses.un1_counterlt13_0_cascade_\
        );

    \I__843\ : InMux
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4164\,
            I => \N__4158\
        );

    \I__841\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4155\
        );

    \I__840\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4152\
        );

    \I__839\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4149\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__4158\,
            I => \arses.counterZ0Z_0\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4155\,
            I => \arses.counterZ0Z_0\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4152\,
            I => \arses.counterZ0Z_0\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4149\,
            I => \arses.counterZ0Z_0\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__833\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4129\
        );

    \I__831\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4126\
        );

    \I__830\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4123\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__4129\,
            I => \N__4118\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4118\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4123\,
            I => \arses.counterZ0Z_1\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__4118\,
            I => \arses.counterZ0Z_1\
        );

    \I__825\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4109\
        );

    \I__824\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4109\,
            I => \arses.counterZ0Z_2\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4106\,
            I => \arses.counterZ0Z_2\
        );

    \I__821\ : InMux
    port map (
            O => \N__4101\,
            I => \arses.un2_counter_cry_1\
        );

    \I__820\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4095\,
            I => \dig1.N_38\
        );

    \I__818\ : InMux
    port map (
            O => \N__4092\,
            I => \N__4089\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4089\,
            I => \dig1.N_35\
        );

    \I__816\ : IoInMux
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4083\,
            I => \N__4080\
        );

    \I__814\ : IoSpan4Mux
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__813\ : Sp12to4
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__812\ : Span12Mux_s6_v
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__811\ : Span12Mux_h
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__810\ : Odrv12
    port map (
            O => \N__4068\,
            I => leds_1_i_0_3
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__4065\,
            I => \N__4061\
        );

    \I__808\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4053\
        );

    \I__807\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4053\
        );

    \I__806\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4053\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4053\,
            I => \dig1.un1_leds114_0\
        );

    \I__804\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4047\,
            I => \dig1.leds_cnst_2\
        );

    \I__802\ : IoInMux
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__800\ : Span4Mux_s1_v
    port map (
            O => \N__4038\,
            I => \N__4035\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__798\ : Sp12to4
    port map (
            O => \N__4032\,
            I => \N__4029\
        );

    \I__797\ : Span12Mux_h
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__796\ : Span12Mux_v
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__795\ : Odrv12
    port map (
            O => \N__4023\,
            I => leds_1_i_0_2
        );

    \I__794\ : IoInMux
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4017\,
            I => \N__4014\
        );

    \I__792\ : Span4Mux_s3_v
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__4011\,
            I => \N__4008\
        );

    \I__790\ : Sp12to4
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__789\ : Span12Mux_s10_h
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4002\,
            I => lcol1_c
        );

    \I__787\ : IoInMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__785\ : Span4Mux_s3_v
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__783\ : Span12Mux_h
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__782\ : Span12Mux_v
    port map (
            O => \N__3984\,
            I => \N__3981\
        );

    \I__781\ : Odrv12
    port map (
            O => \N__3981\,
            I => lcol2_c
        );

    \I__780\ : IoInMux
    port map (
            O => \N__3978\,
            I => \N__3975\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3975\,
            I => \N__3972\
        );

    \I__778\ : Span4Mux_s3_v
    port map (
            O => \N__3972\,
            I => \N__3969\
        );

    \I__777\ : Span4Mux_h
    port map (
            O => \N__3969\,
            I => \N__3966\
        );

    \I__776\ : Span4Mux_v
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__3960\,
            I => \N__3957\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__3957\,
            I => lcol3_c
        );

    \I__772\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3950\
        );

    \I__771\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3943\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3950\,
            I => \N__3940\
        );

    \I__769\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3935\
        );

    \I__768\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3935\
        );

    \I__767\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3930\
        );

    \I__766\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3927\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3943\,
            I => \N__3924\
        );

    \I__764\ : Span4Mux_v
    port map (
            O => \N__3940\,
            I => \N__3919\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3935\,
            I => \N__3919\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__3934\,
            I => \N__3902\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__3933\,
            I => \N__3895\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3930\,
            I => \N__3890\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3927\,
            I => \N__3890\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__3924\,
            I => \N__3885\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__3919\,
            I => \N__3885\
        );

    \I__756\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3882\
        );

    \I__755\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3875\
        );

    \I__754\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3875\
        );

    \I__753\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3875\
        );

    \I__752\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3872\
        );

    \I__751\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3861\
        );

    \I__750\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3861\
        );

    \I__749\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3861\
        );

    \I__748\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3861\
        );

    \I__747\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3861\
        );

    \I__746\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3856\
        );

    \I__745\ : InMux
    port map (
            O => \N__3907\,
            I => \N__3856\
        );

    \I__744\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3849\
        );

    \I__743\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3849\
        );

    \I__742\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3849\
        );

    \I__741\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3844\
        );

    \I__740\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3844\
        );

    \I__739\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3837\
        );

    \I__738\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3837\
        );

    \I__737\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3837\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__3890\,
            I => \colZ0Z_1\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3885\,
            I => \colZ0Z_1\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3882\,
            I => \colZ0Z_1\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3875\,
            I => \colZ0Z_1\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3872\,
            I => \colZ0Z_1\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3861\,
            I => \colZ0Z_1\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3856\,
            I => \colZ0Z_1\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3849\,
            I => \colZ0Z_1\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3844\,
            I => \colZ0Z_1\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3837\,
            I => \colZ0Z_1\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__725\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3806\
        );

    \I__724\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3798\
        );

    \I__723\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3798\
        );

    \I__722\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3795\
        );

    \I__721\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3789\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3806\,
            I => \N__3786\
        );

    \I__719\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3783\
        );

    \I__718\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3778\
        );

    \I__717\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3778\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3798\,
            I => \N__3773\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3795\,
            I => \N__3773\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__3794\,
            I => \N__3770\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__3793\,
            I => \N__3760\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__3792\,
            I => \N__3757\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3789\,
            I => \N__3744\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__3786\,
            I => \N__3735\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3783\,
            I => \N__3735\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3735\
        );

    \I__707\ : Span4Mux_v
    port map (
            O => \N__3773\,
            I => \N__3735\
        );

    \I__706\ : InMux
    port map (
            O => \N__3770\,
            I => \N__3732\
        );

    \I__705\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3729\
        );

    \I__704\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3722\
        );

    \I__703\ : InMux
    port map (
            O => \N__3767\,
            I => \N__3722\
        );

    \I__702\ : InMux
    port map (
            O => \N__3766\,
            I => \N__3722\
        );

    \I__701\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3719\
        );

    \I__700\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3714\
        );

    \I__699\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3714\
        );

    \I__698\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3709\
        );

    \I__697\ : InMux
    port map (
            O => \N__3757\,
            I => \N__3709\
        );

    \I__696\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3704\
        );

    \I__695\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3704\
        );

    \I__694\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3697\
        );

    \I__693\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3697\
        );

    \I__692\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3697\
        );

    \I__691\ : InMux
    port map (
            O => \N__3751\,
            I => \N__3692\
        );

    \I__690\ : InMux
    port map (
            O => \N__3750\,
            I => \N__3692\
        );

    \I__689\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3685\
        );

    \I__688\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3685\
        );

    \I__687\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3685\
        );

    \I__686\ : Odrv4
    port map (
            O => \N__3744\,
            I => \colZ0Z_0\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__3735\,
            I => \colZ0Z_0\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3732\,
            I => \colZ0Z_0\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3729\,
            I => \colZ0Z_0\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3722\,
            I => \colZ0Z_0\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3719\,
            I => \colZ0Z_0\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3714\,
            I => \colZ0Z_0\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3709\,
            I => \colZ0Z_0\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3704\,
            I => \colZ0Z_0\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3697\,
            I => \colZ0Z_0\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3692\,
            I => \colZ0Z_0\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3685\,
            I => \colZ0Z_0\
        );

    \I__674\ : IoInMux
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3657\,
            I => \N__3654\
        );

    \I__672\ : IoSpan4Mux
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__671\ : Span4Mux_s1_v
    port map (
            O => \N__3651\,
            I => \N__3648\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__3648\,
            I => \N__3645\
        );

    \I__669\ : Span12Mux_v
    port map (
            O => \N__3645\,
            I => \N__3642\
        );

    \I__668\ : Span12Mux_h
    port map (
            O => \N__3642\,
            I => \N__3639\
        );

    \I__667\ : Odrv12
    port map (
            O => \N__3639\,
            I => lcol4_c
        );

    \I__666\ : CEMux
    port map (
            O => \N__3636\,
            I => \N__3633\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3633\,
            I => \N__3630\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__3630\,
            I => \N__3624\
        );

    \I__663\ : CEMux
    port map (
            O => \N__3629\,
            I => \N__3621\
        );

    \I__662\ : CEMux
    port map (
            O => \N__3628\,
            I => \N__3618\
        );

    \I__661\ : CEMux
    port map (
            O => \N__3627\,
            I => \N__3615\
        );

    \I__660\ : Span4Mux_v
    port map (
            O => \N__3624\,
            I => \N__3608\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3621\,
            I => \N__3608\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3618\,
            I => \N__3605\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3615\,
            I => \N__3602\
        );

    \I__656\ : CEMux
    port map (
            O => \N__3614\,
            I => \N__3599\
        );

    \I__655\ : CEMux
    port map (
            O => \N__3613\,
            I => \N__3596\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__3608\,
            I => \N__3593\
        );

    \I__653\ : Span4Mux_v
    port map (
            O => \N__3605\,
            I => \N__3586\
        );

    \I__652\ : Span4Mux_v
    port map (
            O => \N__3602\,
            I => \N__3586\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3586\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3596\,
            I => \N__3577\
        );

    \I__649\ : Span4Mux_h
    port map (
            O => \N__3593\,
            I => \N__3574\
        );

    \I__648\ : Span4Mux_v
    port map (
            O => \N__3586\,
            I => \N__3571\
        );

    \I__647\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3564\
        );

    \I__646\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3564\
        );

    \I__645\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3564\
        );

    \I__644\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3559\
        );

    \I__643\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3559\
        );

    \I__642\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3556\
        );

    \I__641\ : Odrv12
    port map (
            O => \N__3577\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__3574\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__639\ : Odrv4
    port map (
            O => \N__3571\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3564\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3559\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3556\,
            I => \clock_out_RNIR6ER_0\
        );

    \I__635\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3540\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3540\,
            I => \N__3537\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__3537\,
            I => \N__3534\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3534\,
            I => \delayConstant_fastZ0Z_2\
        );

    \I__631\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3528\,
            I => \N__3525\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__628\ : Odrv4
    port map (
            O => \N__3522\,
            I => \delayConstant_fastZ0Z_0\
        );

    \I__627\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3516\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3516\,
            I => \dig1.i2_mux\
        );

    \I__625\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3510\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3510\,
            I => \dig1.m23_bm\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__3507\,
            I => \dig1.m29_bm_cascade_\
        );

    \I__622\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3501\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3501\,
            I => \dig1.m23_am\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__3498\,
            I => \dig1.m29_am_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3492\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3492\,
            I => \dig1.m30_ns_1\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__3489\,
            I => \N__3480\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__3488\,
            I => \N__3477\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__3487\,
            I => \N__3474\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__3486\,
            I => \N__3471\
        );

    \I__613\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3462\
        );

    \I__612\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3459\
        );

    \I__611\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3449\
        );

    \I__610\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3449\
        );

    \I__609\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3449\
        );

    \I__608\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3449\
        );

    \I__607\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3444\
        );

    \I__606\ : InMux
    port map (
            O => \N__3470\,
            I => \N__3444\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__3469\,
            I => \N__3441\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__3468\,
            I => \N__3437\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3467\,
            I => \N__3434\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__3466\,
            I => \N__3431\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__3465\,
            I => \N__3428\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3462\,
            I => \N__3425\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3459\,
            I => \N__3422\
        );

    \I__598\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3419\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3449\,
            I => \N__3416\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3444\,
            I => \N__3413\
        );

    \I__595\ : InMux
    port map (
            O => \N__3441\,
            I => \N__3410\
        );

    \I__594\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3403\
        );

    \I__593\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3403\
        );

    \I__592\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3403\
        );

    \I__591\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3398\
        );

    \I__590\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3398\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__3425\,
            I => \delayConstantZ0Z_0\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__3422\,
            I => \delayConstantZ0Z_0\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3419\,
            I => \delayConstantZ0Z_0\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__3416\,
            I => \delayConstantZ0Z_0\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__3413\,
            I => \delayConstantZ0Z_0\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3410\,
            I => \delayConstantZ0Z_0\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3403\,
            I => \delayConstantZ0Z_0\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3398\,
            I => \delayConstantZ0Z_0\
        );

    \I__581\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3375\
        );

    \I__580\ : InMux
    port map (
            O => \N__3380\,
            I => \N__3364\
        );

    \I__579\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3364\
        );

    \I__578\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3364\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3375\,
            I => \N__3361\
        );

    \I__576\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3354\
        );

    \I__575\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3354\
        );

    \I__574\ : InMux
    port map (
            O => \N__3372\,
            I => \N__3354\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__3371\,
            I => \N__3351\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3364\,
            I => \N__3348\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__3361\,
            I => \N__3343\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3354\,
            I => \N__3343\
        );

    \I__569\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3340\
        );

    \I__568\ : Odrv12
    port map (
            O => \N__3348\,
            I => \delayConstantZ0Z_2\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__3343\,
            I => \delayConstantZ0Z_2\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3340\,
            I => \delayConstantZ0Z_2\
        );

    \I__565\ : InMux
    port map (
            O => \N__3333\,
            I => \N__3330\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3330\,
            I => \N__3327\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__3327\,
            I => \dig1.leds_cnst_1\
        );

    \I__562\ : IoInMux
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3321\,
            I => \N__3318\
        );

    \I__560\ : Span4Mux_s3_v
    port map (
            O => \N__3318\,
            I => \N__3315\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__3315\,
            I => \N__3312\
        );

    \I__558\ : Sp12to4
    port map (
            O => \N__3312\,
            I => \N__3309\
        );

    \I__557\ : Span12Mux_s10_h
    port map (
            O => \N__3309\,
            I => \N__3306\
        );

    \I__556\ : Odrv12
    port map (
            O => \N__3306\,
            I => leds_1_i_0_1
        );

    \I__555\ : InMux
    port map (
            O => \N__3303\,
            I => \N__3299\
        );

    \I__554\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3296\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3299\,
            I => \un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3296\,
            I => \un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2\
        );

    \I__551\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3287\
        );

    \I__550\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3284\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3287\,
            I => \un1_delayConstant_cry_3_0_c_RNITFZ0Z062\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3284\,
            I => \un1_delayConstant_cry_3_0_c_RNITFZ0Z062\
        );

    \I__547\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3275\
        );

    \I__546\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3272\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3275\,
            I => \un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3272\,
            I => \un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2\
        );

    \I__543\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3261\
        );

    \I__542\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3261\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3261\,
            I => \un1_delayConstant_cry_1_0_c_RNIP5KDZ0Z2\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__3258\,
            I => \dig1.m8_am_cascade_\
        );

    \I__539\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3252\,
            I => \dig1.m8_bm\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__3249\,
            I => \dig1.N_9_cascade_\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__3246\,
            I => \clock_out_RNIR6ER_0_cascade_\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__3243\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__3240\,
            I => \N__3235\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__3239\,
            I => \N__3232\
        );

    \I__532\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3228\
        );

    \I__531\ : InMux
    port map (
            O => \N__3235\,
            I => \N__3223\
        );

    \I__530\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3223\
        );

    \I__529\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3220\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3228\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3223\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3220\,
            I => \debounceconsolereset.counter_RNINST81Z0Z_4\
        );

    \I__525\ : IoInMux
    port map (
            O => \N__3213\,
            I => \N__3210\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3210\,
            I => \N__3207\
        );

    \I__523\ : Span4Mux_s0_v
    port map (
            O => \N__3207\,
            I => \N__3204\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__3204\,
            I => \N__3198\
        );

    \I__521\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3193\
        );

    \I__520\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3193\
        );

    \I__519\ : InMux
    port map (
            O => \N__3201\,
            I => \N__3189\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__3198\,
            I => \N__3183\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3193\,
            I => \N__3183\
        );

    \I__516\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3180\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3189\,
            I => \N__3177\
        );

    \I__514\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3174\
        );

    \I__513\ : Span4Mux_h
    port map (
            O => \N__3183\,
            I => \N__3171\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3180\,
            I => \N__3168\
        );

    \I__511\ : Span4Mux_v
    port map (
            O => \N__3177\,
            I => \N__3165\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3174\,
            I => \N__3162\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__3171\,
            I => \N__3157\
        );

    \I__508\ : Span4Mux_h
    port map (
            O => \N__3168\,
            I => \N__3157\
        );

    \I__507\ : Sp12to4
    port map (
            O => \N__3165\,
            I => \N__3154\
        );

    \I__506\ : Sp12to4
    port map (
            O => \N__3162\,
            I => \N__3151\
        );

    \I__505\ : Span4Mux_h
    port map (
            O => \N__3157\,
            I => \N__3148\
        );

    \I__504\ : Span12Mux_h
    port map (
            O => \N__3154\,
            I => \N__3145\
        );

    \I__503\ : Span12Mux_v
    port map (
            O => \N__3151\,
            I => \N__3142\
        );

    \I__502\ : Sp12to4
    port map (
            O => \N__3148\,
            I => \N__3139\
        );

    \I__501\ : Span12Mux_v
    port map (
            O => \N__3145\,
            I => \N__3136\
        );

    \I__500\ : Span12Mux_h
    port map (
            O => \N__3142\,
            I => \N__3131\
        );

    \I__499\ : Span12Mux_v
    port map (
            O => \N__3139\,
            I => \N__3131\
        );

    \I__498\ : Odrv12
    port map (
            O => \N__3136\,
            I => masterreset_c
        );

    \I__497\ : Odrv12
    port map (
            O => \N__3131\,
            I => masterreset_c
        );

    \I__496\ : InMux
    port map (
            O => \N__3126\,
            I => \N__3117\
        );

    \I__495\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3117\
        );

    \I__494\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3117\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3117\,
            I => \N__3113\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__3116\,
            I => \N__3110\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__3113\,
            I => \N__3106\
        );

    \I__490\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3101\
        );

    \I__489\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3101\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__3106\,
            I => slowclk
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3101\,
            I => slowclk
        );

    \I__486\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3091\
        );

    \I__485\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3086\
        );

    \I__484\ : InMux
    port map (
            O => \N__3094\,
            I => \N__3086\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3091\,
            I => debouncedn_counter_4
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3086\,
            I => debouncedn_counter_4
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__480\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3073\
        );

    \I__479\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3068\
        );

    \I__478\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3068\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3073\,
            I => debouncedn_counter_1
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3068\,
            I => debouncedn_counter_1
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__3063\,
            I => \N__3058\
        );

    \I__474\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3054\
        );

    \I__473\ : InMux
    port map (
            O => \N__3061\,
            I => \N__3047\
        );

    \I__472\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3047\
        );

    \I__471\ : InMux
    port map (
            O => \N__3057\,
            I => \N__3047\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3054\,
            I => debouncedn_counter_0
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3047\,
            I => debouncedn_counter_0
        );

    \I__468\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3036\
        );

    \I__467\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3033\
        );

    \I__466\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3028\
        );

    \I__465\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3028\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3036\,
            I => \N__3025\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3033\,
            I => debouncedn_counter_2
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3028\,
            I => debouncedn_counter_2
        );

    \I__461\ : Odrv4
    port map (
            O => \N__3025\,
            I => debouncedn_counter_2
        );

    \I__460\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3015\,
            I => \debouncedn.out_cnvZ0Z_1\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3012\,
            I => \N__3008\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3011\,
            I => \N__3005\
        );

    \I__456\ : InMux
    port map (
            O => \N__3008\,
            I => \N__3001\
        );

    \I__455\ : InMux
    port map (
            O => \N__3005\,
            I => \N__2995\
        );

    \I__454\ : InMux
    port map (
            O => \N__3004\,
            I => \N__2995\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3001\,
            I => \N__2992\
        );

    \I__452\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2989\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2995\,
            I => debouncedn_counter_3
        );

    \I__450\ : Odrv4
    port map (
            O => \N__2992\,
            I => debouncedn_counter_3
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2989\,
            I => debouncedn_counter_3
        );

    \I__448\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2979\,
            I => \N__2976\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__2976\,
            I => \N__2973\
        );

    \I__445\ : Sp12to4
    port map (
            O => \N__2973\,
            I => \N__2970\
        );

    \I__444\ : Span12Mux_h
    port map (
            O => \N__2970\,
            I => \N__2967\
        );

    \I__443\ : Span12Mux_v
    port map (
            O => \N__2967\,
            I => \N__2964\
        );

    \I__442\ : Odrv12
    port map (
            O => \N__2964\,
            I => consolereset_c
        );

    \I__441\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2958\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__439\ : Span4Mux_h
    port map (
            O => \N__2955\,
            I => \N__2952\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__2952\,
            I => \N__2949\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__436\ : Span12Mux_h
    port map (
            O => \N__2946\,
            I => \N__2943\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__2943\,
            I => altreset_c
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__2940\,
            I => \out_cnv_cascade_\
        );

    \I__433\ : CascadeMux
    port map (
            O => \N__2937\,
            I => \col_1_1_cascade_\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__2934\,
            I => \dig1.m34_am_cascade_\
        );

    \I__431\ : InMux
    port map (
            O => \N__2931\,
            I => \N__2928\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2928\,
            I => \dig1.m34_bm\
        );

    \I__429\ : InMux
    port map (
            O => \N__2925\,
            I => \debounceconsolereset.un3_counter_cry_1\
        );

    \I__428\ : InMux
    port map (
            O => \N__2922\,
            I => \debounceconsolereset.un3_counter_cry_2\
        );

    \I__427\ : InMux
    port map (
            O => \N__2919\,
            I => \debounceconsolereset.un3_counter_cry_3\
        );

    \I__426\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2913\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2913\,
            I => \debounceconsolereset.un3_counter_cry_2_THRU_CO\
        );

    \I__424\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2907\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2907\,
            I => \debounceconsolereset.un3_counter_cry_1_THRU_CO\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__2904\,
            I => \N__2900\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__2903\,
            I => \N__2897\
        );

    \I__420\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2894\
        );

    \I__419\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2890\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2894\,
            I => \N__2887\
        );

    \I__417\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2882\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2890\,
            I => \N__2876\
        );

    \I__415\ : Span4Mux_h
    port map (
            O => \N__2887\,
            I => \N__2873\
        );

    \I__414\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2870\
        );

    \I__413\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2867\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2882\,
            I => \N__2864\
        );

    \I__411\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2859\
        );

    \I__410\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2859\
        );

    \I__409\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2856\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__2876\,
            I => \delayConstantZ0Z_6\
        );

    \I__407\ : Odrv4
    port map (
            O => \N__2873\,
            I => \delayConstantZ0Z_6\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2870\,
            I => \delayConstantZ0Z_6\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2867\,
            I => \delayConstantZ0Z_6\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__2864\,
            I => \delayConstantZ0Z_6\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2859\,
            I => \delayConstantZ0Z_6\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2856\,
            I => \delayConstantZ0Z_6\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__2841\,
            I => \dig2.m8_am_0_cascade_\
        );

    \I__400\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2835\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2835\,
            I => \dig2.N_9\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__2832\,
            I => \slowclk_0_cascade_\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__396\ : InMux
    port map (
            O => \N__2826\,
            I => \N__2823\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2823\,
            I => slowclk_0
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2820\,
            I => \N__2811\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__2819\,
            I => \N__2808\
        );

    \I__392\ : CascadeMux
    port map (
            O => \N__2818\,
            I => \N__2803\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__2817\,
            I => \N__2800\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__2816\,
            I => \N__2797\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__2815\,
            I => \N__2793\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__2814\,
            I => \N__2790\
        );

    \I__387\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2784\
        );

    \I__386\ : InMux
    port map (
            O => \N__2808\,
            I => \N__2784\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__2807\,
            I => \N__2781\
        );

    \I__384\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2775\
        );

    \I__383\ : InMux
    port map (
            O => \N__2803\,
            I => \N__2775\
        );

    \I__382\ : InMux
    port map (
            O => \N__2800\,
            I => \N__2772\
        );

    \I__381\ : InMux
    port map (
            O => \N__2797\,
            I => \N__2761\
        );

    \I__380\ : InMux
    port map (
            O => \N__2796\,
            I => \N__2761\
        );

    \I__379\ : InMux
    port map (
            O => \N__2793\,
            I => \N__2761\
        );

    \I__378\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2761\
        );

    \I__377\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2761\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2784\,
            I => \N__2758\
        );

    \I__375\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2753\
        );

    \I__374\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2753\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2775\,
            I => \delayConstantZ0Z_4\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2772\,
            I => \delayConstantZ0Z_4\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2761\,
            I => \delayConstantZ0Z_4\
        );

    \I__370\ : Odrv4
    port map (
            O => \N__2758\,
            I => \delayConstantZ0Z_4\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2753\,
            I => \delayConstantZ0Z_4\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__2742\,
            I => \N__2735\
        );

    \I__367\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2724\
        );

    \I__366\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2724\
        );

    \I__365\ : InMux
    port map (
            O => \N__2739\,
            I => \N__2719\
        );

    \I__364\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2719\
        );

    \I__363\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2716\
        );

    \I__362\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2711\
        );

    \I__361\ : InMux
    port map (
            O => \N__2733\,
            I => \N__2711\
        );

    \I__360\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2706\
        );

    \I__359\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2706\
        );

    \I__358\ : InMux
    port map (
            O => \N__2730\,
            I => \N__2701\
        );

    \I__357\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2701\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2724\,
            I => \N__2696\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2719\,
            I => \N__2696\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2716\,
            I => \delayConstantZ0Z_5\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2711\,
            I => \delayConstantZ0Z_5\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2706\,
            I => \delayConstantZ0Z_5\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2701\,
            I => \delayConstantZ0Z_5\
        );

    \I__350\ : Odrv4
    port map (
            O => \N__2696\,
            I => \delayConstantZ0Z_5\
        );

    \I__349\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2682\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2682\,
            I => \dig2.m8_bm_0\
        );

    \I__347\ : InMux
    port map (
            O => \N__2679\,
            I => \N__2675\
        );

    \I__346\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2672\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2675\,
            I => col_1_1
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2672\,
            I => col_1_1
        );

    \I__343\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2664\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2664\,
            I => \olddn_RNISQ7L1Z0Z_0\
        );

    \I__341\ : InMux
    port map (
            O => \N__2661\,
            I => \un1_delayConstant_cry_1\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__2658\,
            I => \N__2655\
        );

    \I__339\ : InMux
    port map (
            O => \N__2655\,
            I => \N__2652\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2652\,
            I => \olddn_RNISQ7L1Z0Z_3\
        );

    \I__337\ : InMux
    port map (
            O => \N__2649\,
            I => \un1_delayConstant_cry_2\
        );

    \I__336\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2643\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2643\,
            I => \olddn_RNISQ7L1Z0Z_1\
        );

    \I__334\ : InMux
    port map (
            O => \N__2640\,
            I => \un1_delayConstant_cry_3\
        );

    \I__333\ : InMux
    port map (
            O => \N__2637\,
            I => \N__2634\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2634\,
            I => \olddn_RNISQ7LZ0Z1\
        );

    \I__331\ : InMux
    port map (
            O => \N__2631\,
            I => \un1_delayConstant_cry_4\
        );

    \I__330\ : InMux
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2625\,
            I => \olddn_RNISQ7L1Z0Z_4\
        );

    \I__328\ : InMux
    port map (
            O => \N__2622\,
            I => \un1_delayConstant_cry_5\
        );

    \I__327\ : InMux
    port map (
            O => \N__2619\,
            I => \un1_delayConstant_cry_6\
        );

    \I__326\ : InMux
    port map (
            O => \N__2616\,
            I => \N__2608\
        );

    \I__325\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2605\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2614\,
            I => \N__2601\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__2613\,
            I => \N__2598\
        );

    \I__322\ : CascadeMux
    port map (
            O => \N__2612\,
            I => \N__2595\
        );

    \I__321\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2590\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2608\,
            I => \N__2585\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2605\,
            I => \N__2585\
        );

    \I__318\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2582\
        );

    \I__317\ : InMux
    port map (
            O => \N__2601\,
            I => \N__2571\
        );

    \I__316\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2571\
        );

    \I__315\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2571\
        );

    \I__314\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2571\
        );

    \I__313\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2571\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2590\,
            I => \delayConstant16_i\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__2585\,
            I => \delayConstant16_i\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2582\,
            I => \delayConstant16_i\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2571\,
            I => \delayConstant16_i\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__2562\,
            I => \N__2557\
        );

    \I__307\ : InMux
    port map (
            O => \N__2561\,
            I => \N__2554\
        );

    \I__306\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2544\
        );

    \I__305\ : InMux
    port map (
            O => \N__2557\,
            I => \N__2541\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2554\,
            I => \N__2538\
        );

    \I__303\ : InMux
    port map (
            O => \N__2553\,
            I => \N__2535\
        );

    \I__302\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2522\
        );

    \I__301\ : InMux
    port map (
            O => \N__2551\,
            I => \N__2522\
        );

    \I__300\ : InMux
    port map (
            O => \N__2550\,
            I => \N__2522\
        );

    \I__299\ : InMux
    port map (
            O => \N__2549\,
            I => \N__2522\
        );

    \I__298\ : InMux
    port map (
            O => \N__2548\,
            I => \N__2522\
        );

    \I__297\ : InMux
    port map (
            O => \N__2547\,
            I => \N__2522\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2544\,
            I => \olddn_RNI1J1RZ0\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2541\,
            I => \olddn_RNI1J1RZ0\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2538\,
            I => \olddn_RNI1J1RZ0\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2535\,
            I => \olddn_RNI1J1RZ0\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2522\,
            I => \olddn_RNI1J1RZ0\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2511\,
            I => \delayConstant16_i_cascade_\
        );

    \I__290\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2505\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2505\,
            I => \oldupZ0\
        );

    \I__288\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2499\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2499\,
            I => \un1_delayConstant_cry_0_c_RNOZ0\
        );

    \I__286\ : CascadeMux
    port map (
            O => \N__2496\,
            I => \N__2493\
        );

    \I__285\ : InMux
    port map (
            O => \N__2493\,
            I => \N__2490\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2490\,
            I => \olddn_RNISQ7L1Z0Z_2\
        );

    \I__283\ : InMux
    port map (
            O => \N__2487\,
            I => \un1_delayConstant_cry_0\
        );

    \I__282\ : InMux
    port map (
            O => \N__2484\,
            I => \N__2481\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2481\,
            I => \dig2.m23_am_0\
        );

    \I__280\ : InMux
    port map (
            O => \N__2478\,
            I => \N__2475\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2475\,
            I => \dig2.m29_am_0\
        );

    \I__278\ : InMux
    port map (
            O => \N__2472\,
            I => \N__2469\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2469\,
            I => \dig2.N_38\
        );

    \I__276\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2463\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2463\,
            I => \dig2.m23_bm_0\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2460\,
            I => \dig2.m34_am_0_cascade_\
        );

    \I__273\ : InMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2454\,
            I => \dig2.m34_bm_0\
        );

    \I__271\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2448\,
            I => \dig2.N_35\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__2445\,
            I => \dig2.leds_cnst_2_cascade_\
        );

    \I__268\ : IoInMux
    port map (
            O => \N__2442\,
            I => \N__2439\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2439\,
            I => \N__2436\
        );

    \I__266\ : Span12Mux_s7_v
    port map (
            O => \N__2436\,
            I => \N__2433\
        );

    \I__265\ : Span12Mux_v
    port map (
            O => \N__2433\,
            I => \N__2430\
        );

    \I__264\ : Span12Mux_h
    port map (
            O => \N__2430\,
            I => \N__2427\
        );

    \I__263\ : Odrv12
    port map (
            O => \N__2427\,
            I => leds_1_i_2
        );

    \I__262\ : InMux
    port map (
            O => \N__2424\,
            I => \N__2421\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2421\,
            I => \olddnZ0\
        );

    \I__260\ : InMux
    port map (
            O => \N__2418\,
            I => \N__2412\
        );

    \I__259\ : InMux
    port map (
            O => \N__2417\,
            I => \N__2412\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2412\,
            I => debounceddn
        );

    \I__257\ : InMux
    port map (
            O => \N__2409\,
            I => \N__2404\
        );

    \I__256\ : InMux
    port map (
            O => \N__2408\,
            I => \N__2399\
        );

    \I__255\ : InMux
    port map (
            O => \N__2407\,
            I => \N__2399\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2404\,
            I => \dig2.un1_leds114_0\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2399\,
            I => \dig2.un1_leds114_0\
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2394\,
            I => \dig2.i2_mux_cascade_\
        );

    \I__251\ : InMux
    port map (
            O => \N__2391\,
            I => \N__2388\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2388\,
            I => \dig2.leds_cnst_1\
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__2385\,
            I => \dig2.m29_bm_0_cascade_\
        );

    \I__248\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2379\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2379\,
            I => \dig2.m30_ns_1\
        );

    \I__246\ : IoInMux
    port map (
            O => \N__2376\,
            I => \N__2373\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2373\,
            I => \N__2370\
        );

    \I__244\ : IoSpan4Mux
    port map (
            O => \N__2370\,
            I => \N__2367\
        );

    \I__243\ : Span4Mux_s2_v
    port map (
            O => \N__2367\,
            I => \N__2364\
        );

    \I__242\ : Sp12to4
    port map (
            O => \N__2364\,
            I => \N__2361\
        );

    \I__241\ : Span12Mux_s10_v
    port map (
            O => \N__2361\,
            I => \N__2358\
        );

    \I__240\ : Span12Mux_v
    port map (
            O => \N__2358\,
            I => \N__2355\
        );

    \I__239\ : Span12Mux_h
    port map (
            O => \N__2355\,
            I => \N__2352\
        );

    \I__238\ : Odrv12
    port map (
            O => \N__2352\,
            I => \arse.divseven.io_0_D_IN_0\
        );

    \I__237\ : IoInMux
    port map (
            O => \N__2349\,
            I => \N__2346\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2346\,
            I => \N__2343\
        );

    \I__235\ : Span12Mux_s8_h
    port map (
            O => \N__2343\,
            I => \N__2340\
        );

    \I__234\ : Odrv12
    port map (
            O => \N__2340\,
            I => masterreset_c_i
        );

    \I__233\ : IoInMux
    port map (
            O => \N__2337\,
            I => \N__2334\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2334\,
            I => \N__2331\
        );

    \I__231\ : IoSpan4Mux
    port map (
            O => \N__2331\,
            I => \N__2328\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__2328\,
            I => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\
        );

    \I__229\ : InMux
    port map (
            O => \N__2325\,
            I => \N__2322\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2322\,
            I => \N__2319\
        );

    \I__227\ : Span4Mux_v
    port map (
            O => \N__2319\,
            I => \N__2316\
        );

    \I__226\ : Sp12to4
    port map (
            O => \N__2316\,
            I => \N__2313\
        );

    \I__225\ : Span12Mux_h
    port map (
            O => \N__2313\,
            I => \N__2310\
        );

    \I__224\ : Span12Mux_v
    port map (
            O => \N__2310\,
            I => \N__2307\
        );

    \I__223\ : Odrv12
    port map (
            O => \N__2307\,
            I => deldn_c
        );

    \I__222\ : IoInMux
    port map (
            O => \N__2304\,
            I => \N__2301\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2301\,
            I => \N__2298\
        );

    \I__220\ : Span4Mux_s0_v
    port map (
            O => \N__2298\,
            I => \N__2295\
        );

    \I__219\ : Sp12to4
    port map (
            O => \N__2295\,
            I => \N__2292\
        );

    \I__218\ : Span12Mux_h
    port map (
            O => \N__2292\,
            I => \N__2289\
        );

    \I__217\ : Span12Mux_v
    port map (
            O => \N__2289\,
            I => \N__2286\
        );

    \I__216\ : Odrv12
    port map (
            O => \N__2286\,
            I => leds_1_i_1
        );

    \I__215\ : IoInMux
    port map (
            O => \N__2283\,
            I => \N__2280\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2280\,
            I => \N__2277\
        );

    \I__213\ : Span4Mux_s3_v
    port map (
            O => \N__2277\,
            I => \N__2274\
        );

    \I__212\ : Span4Mux_v
    port map (
            O => \N__2274\,
            I => \N__2271\
        );

    \I__211\ : Sp12to4
    port map (
            O => \N__2271\,
            I => \N__2268\
        );

    \I__210\ : Span12Mux_h
    port map (
            O => \N__2268\,
            I => \N__2265\
        );

    \I__209\ : Span12Mux_v
    port map (
            O => \N__2265\,
            I => \N__2262\
        );

    \I__208\ : Odrv12
    port map (
            O => \N__2262\,
            I => leds_1_i_3
        );

    \I__207\ : ClkMux
    port map (
            O => \N__2259\,
            I => \N__2256\
        );

    \I__206\ : GlobalMux
    port map (
            O => \N__2256\,
            I => \N__2253\
        );

    \I__205\ : gio2CtrlBuf
    port map (
            O => \N__2253\,
            I => \arse.un1_io_0_1_g\
        );

    \I__204\ : IoInMux
    port map (
            O => \N__2250\,
            I => \N__2247\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__2247\,
            I => \N__2244\
        );

    \I__202\ : Span4Mux_s1_v
    port map (
            O => \N__2244\,
            I => \N__2241\
        );

    \I__201\ : Sp12to4
    port map (
            O => \N__2241\,
            I => \N__2238\
        );

    \I__200\ : Span12Mux_h
    port map (
            O => \N__2238\,
            I => \N__2235\
        );

    \I__199\ : Span12Mux_v
    port map (
            O => \N__2235\,
            I => \N__2232\
        );

    \I__198\ : Span12Mux_v
    port map (
            O => \N__2232\,
            I => \N__2229\
        );

    \I__197\ : Odrv12
    port map (
            O => \N__2229\,
            I => \top_pll_nrtthrth.PLLOUTCORE\
        );

    \INVarse.diveight.dout_0C\ : INV
    port map (
            O => \INVarse.diveight.dout_0C_net\,
            I => \N__5397\
        );

    \INVarse.apusynclatchedC\ : INV
    port map (
            O => \INVarse.apusynclatchedC_net\,
            I => \N__2259\
        );

    \INVarse.cpuclkresetC\ : INV
    port map (
            O => \INVarse.cpuclkresetC_net\,
            I => \N__5393\
        );

    \INVarse.divseven.dout_0C\ : INV
    port map (
            O => \INVarse.divseven.dout_0C_net\,
            I => \N__5392\
        );

    \INVarse.cpuresetcount_0C\ : INV
    port map (
            O => \INVarse.cpuresetcount_0C_net\,
            I => \N__5389\
        );

    \INVarse.cpuresetoutregC\ : INV
    port map (
            O => \INVarse.cpuresetoutregC_net\,
            I => \N__5387\
        );

    \INVarse.doingsevenC\ : INV
    port map (
            O => \INVarse.doingsevenC_net\,
            I => \N__5388\
        );

    \IN_MUX_bfv_21_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_11_0_\
        );

    \IN_MUX_bfv_22_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_8_0_\
        );

    \IN_MUX_bfv_23_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_10_0_\
        );

    \IN_MUX_bfv_23_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \arses.un2_counter_cry_8\,
            carryinitout => \bfn_23_11_0_\
        );

    \IN_MUX_bfv_24_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_8_0_\
        );

    \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2250\,
            GLOBALBUFFEROUTPUT => \PLLOUTCORE_g\
        );

    \arse.divseven.io_0_RNIIG08\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2376\,
            GLOBALBUFFEROUTPUT => \arse.un1_io_0_1_g\
        );

    \masterreset_ibuf_RNIKP26_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2349\,
            GLOBALBUFFEROUTPUT => masterreset_c_i_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \masterreset_ibuf_RNIKP26_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3188\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => masterreset_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.out_e_0_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => debounceddn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5293\,
            ce => \N__5237\,
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_1_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000011"
        )
    port map (
            in0 => \N__2391\,
            in1 => \N__3953\,
            in2 => \N__3816\,
            in3 => \N__2409\,
            lcout => leds_1_i_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5297\,
            ce => \N__3629\,
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_3_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010001100"
        )
    port map (
            in0 => \N__2472\,
            in1 => \N__2408\,
            in2 => \N__5076\,
            in3 => \N__2451\,
            lcout => leds_1_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5300\,
            ce => \N__3636\,
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m30_ns_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111100"
        )
    port map (
            in0 => \N__2484\,
            in1 => \N__2478\,
            in2 => \N__2904\,
            in3 => \N__2382\,
            lcout => OPEN,
            ltout => \dig2.leds_cnst_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_1_i_2_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2407\,
            in2 => \N__2445\,
            in3 => \N__3809\,
            lcout => leds_1_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5300\,
            ce => \N__3636\,
            sr => \_gnd_net_\
        );

    \olddn_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2418\,
            lcout => \olddnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNI1J1R_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2424\,
            in2 => \_gnd_net_\,
            in3 => \N__2417\,
            lcout => \olddn_RNI1J1RZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNISQ7L1_3_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2604\,
            in2 => \_gnd_net_\,
            in3 => \N__2553\,
            lcout => \olddn_RNISQ7L1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.un1_leds114_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110111111111"
        )
    port map (
            in0 => \N__2886\,
            in1 => \N__2806\,
            in2 => \N__5070\,
            in3 => \N__2734\,
            lcout => \dig2.un1_leds114_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m11_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110011100011"
        )
    port map (
            in0 => \N__2733\,
            in1 => \N__3918\,
            in2 => \N__2818\,
            in3 => \N__3769\,
            lcout => OPEN,
            ltout => \dig2.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m13_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110111"
        )
    port map (
            in0 => \N__5056\,
            in1 => \N__2885\,
            in2 => \N__2394\,
            in3 => \N__2838\,
            lcout => \dig2.leds_cnst_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m29_bm_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101001011101"
        )
    port map (
            in0 => \N__3766\,
            in1 => \N__2731\,
            in2 => \N__2814\,
            in3 => \N__3910\,
            lcout => OPEN,
            ltout => \dig2.m29_bm_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m30_ns_1_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100100111011"
        )
    port map (
            in0 => \N__2880\,
            in1 => \N__5071\,
            in2 => \N__2385\,
            in3 => \N__2466\,
            lcout => \dig2.m30_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m23_am_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110101101"
        )
    port map (
            in0 => \N__3911\,
            in1 => \N__2730\,
            in2 => \N__3793\,
            in3 => \N__2796\,
            lcout => \dig2.m23_am_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m29_am_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010101"
        )
    port map (
            in0 => \N__3767\,
            in1 => \N__2732\,
            in2 => \N__2815\,
            in3 => \N__3912\,
            lcout => \dig2.m29_am_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m37_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3768\,
            in1 => \N__3913\,
            in2 => \N__2816\,
            in3 => \N__2881\,
            lcout => \dig2.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m23_bm_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000110"
        )
    port map (
            in0 => \N__3909\,
            in1 => \N__2729\,
            in2 => \N__3792\,
            in3 => \N__2789\,
            lcout => \dig2.m23_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m34_bm_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100110111"
        )
    port map (
            in0 => \N__2740\,
            in1 => \N__3914\,
            in2 => \N__2819\,
            in3 => \N__3765\,
            lcout => \dig2.m34_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m34_am_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__2741\,
            in1 => \_gnd_net_\,
            in2 => \N__2820\,
            in3 => \N__2678\,
            lcout => OPEN,
            ltout => \dig2.m34_am_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m34_ns_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2893\,
            in2 => \N__2460\,
            in3 => \N__2457\,
            lcout => \dig2.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_fast_0_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__3484\,
            in1 => \N__2611\,
            in2 => \_gnd_net_\,
            in3 => \N__2560\,
            lcout => \delayConstant_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5295\,
            ce => 'H',
            sr => \N__4444\
        );

    \arses.counter_1_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4132\,
            in1 => \N__4167\,
            in2 => \_gnd_net_\,
            in3 => \N__4557\,
            lcout => \arses.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5295\,
            ce => 'H',
            sr => \N__4444\
        );

    \olddn_RNISQ7L1_0_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2594\,
            in2 => \_gnd_net_\,
            in3 => \N__2549\,
            lcout => \olddn_RNISQ7L1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oldup_RNIR76Q_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__3201\,
            in1 => \N__2508\,
            in2 => \_gnd_net_\,
            in3 => \N__5327\,
            lcout => \delayConstant16_i\,
            ltout => \delayConstant16_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_0_c_RNO_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \N__3485\,
            in1 => \_gnd_net_\,
            in2 => \N__2511\,
            in3 => \N__2547\,
            lcout => \un1_delayConstant_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNISQ7L1_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__2551\,
            in1 => \_gnd_net_\,
            in2 => \N__2613\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNISQ7LZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oldup_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5328\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \oldupZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNISQ7L1_1_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__2550\,
            in1 => \_gnd_net_\,
            in2 => \N__2612\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNISQ7L1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNISQ7L1_2_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2593\,
            in2 => \_gnd_net_\,
            in3 => \N__2548\,
            lcout => \olddn_RNISQ7L1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \olddn_RNISQ7L1_4_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__2552\,
            in1 => \_gnd_net_\,
            in2 => \N__2614\,
            in3 => \_gnd_net_\,
            lcout => \olddn_RNISQ7L1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_0_c_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2502\,
            in2 => \N__3469\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_11_0_\,
            carryout => \un1_delayConstant_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_1_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4979\,
            in2 => \N__2496\,
            in3 => \N__2487\,
            lcout => \delayConstantZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_0\,
            carryout => \un1_delayConstant_cry_1\,
            clk => \N__5301\,
            ce => 'H',
            sr => \N__4442\
        );

    \un1_delayConstant_cry_1_0_c_RNIP5KD2_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2667\,
            in2 => \N__3371\,
            in3 => \N__2661\,
            lcout => \un1_delayConstant_cry_1_0_c_RNIP5KDZ0Z2\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_1\,
            carryout => \un1_delayConstant_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_3_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4795\,
            in2 => \N__2658\,
            in3 => \N__2649\,
            lcout => \delayConstantZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_2\,
            carryout => \un1_delayConstant_cry_3\,
            clk => \N__5301\,
            ce => 'H',
            sr => \N__4442\
        );

    \un1_delayConstant_cry_3_0_c_RNITF062_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2646\,
            in2 => \N__2817\,
            in3 => \N__2640\,
            lcout => \un1_delayConstant_cry_3_0_c_RNITFZ0Z062\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_3\,
            carryout => \un1_delayConstant_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_4_0_c_RNIVK6A2_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2637\,
            in2 => \N__2742\,
            in3 => \N__2631\,
            lcout => \un1_delayConstant_cry_4_0_c_RNIVK6AZ0Z2\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_4\,
            carryout => \un1_delayConstant_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_delayConstant_cry_5_0_c_RNI1QCE2_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2628\,
            in2 => \N__2903\,
            in3 => \N__2622\,
            lcout => \un1_delayConstant_cry_5_0_c_RNI1QCEZ0Z2\,
            ltout => OPEN,
            carryin => \un1_delayConstant_cry_5\,
            carryout => \un1_delayConstant_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_7_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__5060\,
            in1 => \N__2616\,
            in2 => \N__2562\,
            in3 => \N__2619\,
            lcout => \delayConstantZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5301\,
            ce => 'H',
            sr => \N__4442\
        );

    \delayConstant_0_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__3458\,
            in1 => \N__2615\,
            in2 => \_gnd_net_\,
            in3 => \N__2561\,
            lcout => \delayConstantZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5303\,
            ce => 'H',
            sr => \N__4441\
        );

    \delayConstant_5_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3278\,
            lcout => \delayConstantZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5303\,
            ce => 'H',
            sr => \N__4441\
        );

    \delayConstant_4_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3290\,
            lcout => \delayConstantZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5303\,
            ce => 'H',
            sr => \N__4441\
        );

    \delayConstant_6_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3302\,
            lcout => \delayConstantZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5303\,
            ce => 'H',
            sr => \N__4441\
        );

    \dig2.leds_cnst_3_1__m8_am_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000001111010"
        )
    port map (
            in0 => \N__2739\,
            in1 => \N__3898\,
            in2 => \N__2807\,
            in3 => \N__3748\,
            lcout => OPEN,
            ltout => \dig2.m8_am_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m8_ns_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2879\,
            in1 => \_gnd_net_\,
            in2 => \N__2841\,
            in3 => \N__2685\,
            lcout => \dig2.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__3192\,
            in1 => \N__3124\,
            in2 => \_gnd_net_\,
            in3 => \N__4555\,
            lcout => slowclk_0,
            ltout => \slowclk_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \col_0_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__3125\,
            in1 => \_gnd_net_\,
            in2 => \N__2832\,
            in3 => \N__3749\,
            lcout => \colZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \col_1_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__3899\,
            in1 => \N__2679\,
            in2 => \N__2829\,
            in3 => \N__3126\,
            lcout => \colZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig2.leds_cnst_3_1__m8_bm_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3747\,
            in1 => \N__2780\,
            in2 => \N__3933\,
            in3 => \N__2738\,
            lcout => \dig2.m8_bm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m34_bm_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100110111"
        )
    port map (
            in0 => \N__4993\,
            in1 => \N__3908\,
            in2 => \N__3486\,
            in3 => \N__3756\,
            lcout => \dig1.m34_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m11x_i_o2_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3907\,
            in2 => \_gnd_net_\,
            in3 => \N__3755\,
            lcout => col_1_1,
            ltout => \col_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m34_am_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3470\,
            in2 => \N__2937\,
            in3 => \N__4994\,
            lcout => OPEN,
            ltout => \dig1.m34_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m34_ns_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3381\,
            in2 => \N__2934\,
            in3 => \N__2931\,
            lcout => \dig1.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_1_c_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3062\,
            in2 => \N__3081\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_8_0_\,
            carryout => \debounceconsolereset.un3_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_1_THRU_LUT4_0_LC_22_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3039\,
            in2 => \_gnd_net_\,
            in3 => \N__2925\,
            lcout => \debounceconsolereset.un3_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_1\,
            carryout => \debounceconsolereset.un3_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.un3_counter_cry_2_THRU_LUT4_0_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3004\,
            in2 => \_gnd_net_\,
            in3 => \N__2922\,
            lcout => \debounceconsolereset.un3_counter_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \debounceconsolereset.un3_counter_cry_2\,
            carryout => \debounceconsolereset.un3_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_4_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__3096\,
            in1 => \N__3583\,
            in2 => \N__3239\,
            in3 => \N__2919\,
            lcout => debouncedn_counter_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_3_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__2916\,
            in1 => \N__3585\,
            in2 => \N__3011\,
            in3 => \N__3238\,
            lcout => debouncedn_counter_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_2_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__2910\,
            in1 => \N__3584\,
            in2 => \N__3240\,
            in3 => \N__3040\,
            lcout => debouncedn_counter_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_RNIR6ER_0_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__3203\,
            in1 => \N__3109\,
            in2 => \_gnd_net_\,
            in3 => \N__4500\,
            lcout => \clock_out_RNIR6ER_0\,
            ltout => \clock_out_RNIR6ER_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_RNINST81_4_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__3095\,
            in1 => \N__3000\,
            in2 => \N__3246\,
            in3 => \N__3041\,
            lcout => \debounceconsolereset.counter_RNINST81Z0Z_4\,
            ltout => \debounceconsolereset.counter_RNINST81Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_0_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__3061\,
            in1 => \_gnd_net_\,
            in2 => \N__3243\,
            in3 => \N__3581\,
            lcout => debouncedn_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.counter_1_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__3077\,
            in1 => \N__3231\,
            in2 => \N__3063\,
            in3 => \N__3582\,
            lcout => debouncedn_counter_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.clock_out_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__4501\,
            in1 => \_gnd_net_\,
            in2 => \N__3116\,
            in3 => \N__3202\,
            lcout => slowclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.out_cnv_1_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3094\,
            in1 => \N__3076\,
            in2 => \_gnd_net_\,
            in3 => \N__3057\,
            lcout => \debouncedn.out_cnvZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI1L5_2_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4343\,
            in1 => \N__4112\,
            in2 => \_gnd_net_\,
            in3 => \N__4161\,
            lcout => \arses.un1_counterlto4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debouncedn.out_cnv_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__3042\,
            in1 => \N__3018\,
            in2 => \N__3012\,
            in3 => \N__3580\,
            lcout => out_cnv,
            ltout => \out_cnv_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__2982\,
            in1 => \N__2961\,
            in2 => \N__2940\,
            in3 => \N__5524\,
            lcout => debouncedconsolereset,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delayConstant_2_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3266\,
            lcout => \delayConstantZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5304\,
            ce => 'H',
            sr => \N__4443\
        );

    \delayConstant_fast_6_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3303\,
            lcout => \delayConstant_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5304\,
            ce => 'H',
            sr => \N__4443\
        );

    \delayConstant_fast_4_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3291\,
            lcout => \delayConstant_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5304\,
            ce => 'H',
            sr => \N__4443\
        );

    \arses.counter_0_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4163\,
            in2 => \_gnd_net_\,
            in3 => \N__4556\,
            lcout => \arses.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5304\,
            ce => 'H',
            sr => \N__4443\
        );

    \delayConstant_fast_5_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3279\,
            lcout => \delayConstant_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5304\,
            ce => 'H',
            sr => \N__4443\
        );

    \delayConstant_fast_2_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delayConstant_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5304\,
            ce => 'H',
            sr => \N__4443\
        );

    \dig1.leds_cnst_3_1__m23_bm_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110110"
        )
    port map (
            in0 => \N__4960\,
            in1 => \N__3901\,
            in2 => \N__3466\,
            in3 => \N__3750\,
            lcout => \dig1.m23_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m8_bm_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4959\,
            in1 => \N__3900\,
            in2 => \N__3465\,
            in3 => \N__3751\,
            lcout => \dig1.m8_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m8_am_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000001111010"
        )
    port map (
            in0 => \N__4982\,
            in1 => \N__3906\,
            in2 => \N__3468\,
            in3 => \N__3754\,
            lcout => OPEN,
            ltout => \dig1.m8_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m8_ns_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__3373\,
            in1 => \_gnd_net_\,
            in2 => \N__3258\,
            in3 => \N__3255\,
            lcout => OPEN,
            ltout => \dig1.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m13_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110101111"
        )
    port map (
            in0 => \N__4800\,
            in1 => \N__3519\,
            in2 => \N__3249\,
            in3 => \N__3374\,
            lcout => \dig1.leds_cnst_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m11_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010100101"
        )
    port map (
            in0 => \N__3752\,
            in1 => \N__4980\,
            in2 => \N__3934\,
            in3 => \N__3440\,
            lcout => \dig1.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m29_bm_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111010110011"
        )
    port map (
            in0 => \N__4981\,
            in1 => \N__3905\,
            in2 => \N__3467\,
            in3 => \N__3753\,
            lcout => OPEN,
            ltout => \dig1.m29_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m30_ns_1_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__3372\,
            in1 => \N__3513\,
            in2 => \N__3507\,
            in3 => \N__4799\,
            lcout => \dig1.m30_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m23_am_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001111011"
        )
    port map (
            in0 => \N__4995\,
            in1 => \N__3915\,
            in2 => \N__3487\,
            in3 => \N__3763\,
            lcout => \dig1.m23_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.un1_leds114_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111110111"
        )
    port map (
            in0 => \N__4997\,
            in1 => \N__3379\,
            in2 => \N__3489\,
            in3 => \N__4801\,
            lcout => \dig1.un1_leds114_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m29_am_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111111"
        )
    port map (
            in0 => \N__4996\,
            in1 => \N__3916\,
            in2 => \N__3488\,
            in3 => \N__3764\,
            lcout => OPEN,
            ltout => \dig1.m29_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m30_ns_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111010"
        )
    port map (
            in0 => \N__3378\,
            in1 => \N__3504\,
            in2 => \N__3498\,
            in3 => \N__3495\,
            lcout => \dig1.leds_cnst_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_cnst_3_1__m37_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3483\,
            in1 => \N__3917\,
            in2 => \N__3794\,
            in3 => \N__3380\,
            lcout => \dig1.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_1_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010011"
        )
    port map (
            in0 => \N__3333\,
            in1 => \N__3804\,
            in2 => \N__4065\,
            in3 => \N__3947\,
            lcout => leds_1_i_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5309\,
            ce => \N__3614\,
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_3_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001100000000"
        )
    port map (
            in0 => \N__4098\,
            in1 => \N__4092\,
            in2 => \N__4812\,
            in3 => \N__4064\,
            lcout => leds_1_i_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5309\,
            ce => \N__3614\,
            sr => \_gnd_net_\
        );

    \dig1.leds_1_i_2_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__3803\,
            in1 => \N__4060\,
            in2 => \_gnd_net_\,
            in3 => \N__4050\,
            lcout => leds_1_i_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5309\,
            ce => \N__3614\,
            sr => \_gnd_net_\
        );

    \lcolreg_0_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3805\,
            in2 => \_gnd_net_\,
            in3 => \N__3946\,
            lcout => lcol1_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5310\,
            ce => \N__3613\,
            sr => \_gnd_net_\
        );

    \lcolreg_1_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3948\,
            in2 => \_gnd_net_\,
            in3 => \N__3811\,
            lcout => lcol2_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5311\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \lcolreg_2_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3949\,
            in2 => \_gnd_net_\,
            in3 => \N__3812\,
            lcout => lcol3_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5311\,
            ce => \N__3627\,
            sr => \_gnd_net_\
        );

    \lcolreg_3_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3954\,
            in2 => \_gnd_net_\,
            in3 => \N__3810\,
            lcout => lcol4_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5312\,
            ce => \N__3628\,
            sr => \_gnd_net_\
        );

    \arse.doingseven_LC_23_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__5725\,
            in1 => \N__4709\,
            in2 => \_gnd_net_\,
            in3 => \N__4359\,
            lcout => \arse.doingsevenZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.doingsevenC_net\,
            ce => 'H',
            sr => \N__5123\
        );

    \arse.cpuresetoutreg_RNO_6_LC_23_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__3543\,
            in1 => \N__3531\,
            in2 => \N__4674\,
            in3 => \N__4644\,
            lcout => OPEN,
            ltout => \arse.g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_3_LC_23_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4716\,
            in2 => \N__4215\,
            in3 => \N__4830\,
            lcout => OPEN,
            ltout => \arse.g0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_0_LC_23_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5730\,
            in1 => \N__4905\,
            in2 => \N__4212\,
            in3 => \N__4350\,
            lcout => OPEN,
            ltout => \arse.cpuresetoutreg_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4209\,
            in3 => \N__4196\,
            lcout => \arse.cpuresetoutregZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuresetoutregC_net\,
            ce => 'H',
            sr => \N__5124\
        );

    \arses.counter_RNIA58_5_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4283\,
            in1 => \N__4298\,
            in2 => \N__4269\,
            in3 => \N__4313\,
            lcout => OPEN,
            ltout => \arses.un1_counterlto8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOKH_1_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4328\,
            in1 => \N__4133\,
            in2 => \N__4182\,
            in3 => \N__4179\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNI04C4_9_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4611\,
            in1 => \N__4233\,
            in2 => \N__4173\,
            in3 => \N__4251\,
            lcout => OPEN,
            ltout => \arses.un1_counterlt13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_RNIOS0A_14_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__4593\,
            in1 => \N__4464\,
            in2 => \N__4170\,
            in3 => \N__4575\,
            lcout => \arses.counter8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.un2_counter_cry_1_c_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4162\,
            in2 => \N__4140\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_23_10_0_\,
            carryout => \arses.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arses.counter_2_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4551\,
            in1 => \N__4113\,
            in2 => \_gnd_net_\,
            in3 => \N__4101\,
            lcout => \arses.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_1\,
            carryout => \arses.un2_counter_cry_2\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_3_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4533\,
            in1 => \N__4344\,
            in2 => \_gnd_net_\,
            in3 => \N__4332\,
            lcout => \arses.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_2\,
            carryout => \arses.un2_counter_cry_3\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_4_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4552\,
            in1 => \N__4329\,
            in2 => \_gnd_net_\,
            in3 => \N__4317\,
            lcout => \arses.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_3\,
            carryout => \arses.un2_counter_cry_4\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_5_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4534\,
            in1 => \N__4314\,
            in2 => \_gnd_net_\,
            in3 => \N__4302\,
            lcout => \arses.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_4\,
            carryout => \arses.un2_counter_cry_5\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_6_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4553\,
            in1 => \N__4299\,
            in2 => \_gnd_net_\,
            in3 => \N__4287\,
            lcout => \arses.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_5\,
            carryout => \arses.un2_counter_cry_6\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_7_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4535\,
            in1 => \N__4284\,
            in2 => \_gnd_net_\,
            in3 => \N__4272\,
            lcout => \arses.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_6\,
            carryout => \arses.un2_counter_cry_7\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_8_LC_23_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4554\,
            in1 => \N__4268\,
            in2 => \_gnd_net_\,
            in3 => \N__4254\,
            lcout => \arses.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_7\,
            carryout => \arses.un2_counter_cry_8\,
            clk => \N__5305\,
            ce => 'H',
            sr => \N__4446\
        );

    \arses.counter_9_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4547\,
            in1 => \N__4250\,
            in2 => \_gnd_net_\,
            in3 => \N__4236\,
            lcout => \arses.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_23_11_0_\,
            carryout => \arses.un2_counter_cry_9\,
            clk => \N__5307\,
            ce => 'H',
            sr => \N__4445\
        );

    \arses.counter_10_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4548\,
            in1 => \N__4232\,
            in2 => \_gnd_net_\,
            in3 => \N__4218\,
            lcout => \arses.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_9\,
            carryout => \arses.un2_counter_cry_10\,
            clk => \N__5307\,
            ce => 'H',
            sr => \N__4445\
        );

    \arses.counter_11_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4545\,
            in1 => \N__4610\,
            in2 => \_gnd_net_\,
            in3 => \N__4596\,
            lcout => \arses.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_10\,
            carryout => \arses.un2_counter_cry_11\,
            clk => \N__5307\,
            ce => 'H',
            sr => \N__4445\
        );

    \arses.counter_12_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4549\,
            in1 => \N__4592\,
            in2 => \_gnd_net_\,
            in3 => \N__4578\,
            lcout => \arses.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_11\,
            carryout => \arses.un2_counter_cry_12\,
            clk => \N__5307\,
            ce => 'H',
            sr => \N__4445\
        );

    \arses.counter_13_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4546\,
            in1 => \N__4574\,
            in2 => \_gnd_net_\,
            in3 => \N__4560\,
            lcout => \arses.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \arses.un2_counter_cry_12\,
            carryout => \arses.un2_counter_cry_13\,
            clk => \N__5307\,
            ce => 'H',
            sr => \N__4445\
        );

    \arses.counter_14_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4550\,
            in1 => \N__4460\,
            in2 => \_gnd_net_\,
            in3 => \N__4467\,
            lcout => \arses.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5307\,
            ce => 'H',
            sr => \N__4445\
        );

    \CONSTANT_ONE_LUT4_LC_23_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.doingseven_RNO_0_LC_24_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4686\,
            in1 => \N__4647\,
            in2 => \N__4695\,
            in3 => \N__4739\,
            lcout => \arse.doingseven3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_RNIB4QP_0_LC_24_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4668\,
            in2 => \_gnd_net_\,
            in3 => \N__5022\,
            lcout => \arse.doingseven3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_4_LC_24_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__4669\,
            in1 => \N__4759\,
            in2 => \N__5025\,
            in3 => \N__4849\,
            lcout => OPEN,
            ltout => \arse.g0_i_a3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_1_LC_24_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4929\,
            in1 => \N__4870\,
            in2 => \N__4353\,
            in3 => \N__4737\,
            lcout => \arse.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_RNIATKJ1_7_LC_24_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4869\,
            in1 => \N__4758\,
            in2 => \N__4932\,
            in3 => \N__4850\,
            lcout => \arse.doingseven3_6\,
            ltout => \arse.doingseven3_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuclkreset_RNO_0_LC_24_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4685\,
            in1 => \N__4646\,
            in2 => \N__4677\,
            in3 => \N__4738\,
            lcout => \arse.doingseven4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetcount_0_LC_24_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4670\,
            in2 => \N__5729\,
            in3 => \N__5724\,
            lcout => \arse.cpuresetcountZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_24_8_0_\,
            carryout => \arse.un1_cpuresetcount_1_cry_0\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_1_LC_24_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5024\,
            in2 => \_gnd_net_\,
            in3 => \N__4650\,
            lcout => \arse.cpuresetcountZ0Z_1\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_0\,
            carryout => \arse.un1_cpuresetcount_1_cry_1\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_2_LC_24_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4645\,
            in2 => \_gnd_net_\,
            in3 => \N__4626\,
            lcout => \arse.cpuresetcountZ0Z_2\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_1\,
            carryout => \arse.un1_cpuresetcount_1_cry_2\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_3_LC_24_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4740\,
            in2 => \_gnd_net_\,
            in3 => \N__4623\,
            lcout => \arse.cpuresetcountZ0Z_3\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_2\,
            carryout => \arse.un1_cpuresetcount_1_cry_3\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_4_LC_24_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4763\,
            in2 => \_gnd_net_\,
            in3 => \N__4620\,
            lcout => \arse.cpuresetcountZ0Z_4\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_3\,
            carryout => \arse.un1_cpuresetcount_1_cry_4\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_5_LC_24_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4851\,
            in2 => \_gnd_net_\,
            in3 => \N__4617\,
            lcout => \arse.cpuresetcountZ0Z_5\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_4\,
            carryout => \arse.un1_cpuresetcount_1_cry_5\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_6_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4874\,
            in2 => \_gnd_net_\,
            in3 => \N__4614\,
            lcout => \arse.cpuresetcountZ0Z_6\,
            ltout => OPEN,
            carryin => \arse.un1_cpuresetcount_1_cry_5\,
            carryout => \arse.un1_cpuresetcount_1_cry_6\,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetcount_7_LC_24_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4931\,
            in2 => \_gnd_net_\,
            in3 => \N__5079\,
            lcout => \arse.cpuresetcountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuresetcount_0C_net\,
            ce => 'H',
            sr => \N__5115\
        );

    \arse.cpuresetoutreg_RNO_2_LC_24_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__5075\,
            in1 => \N__5023\,
            in2 => \N__5001\,
            in3 => \N__4930\,
            lcout => \arse.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_7_LC_24_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__4899\,
            in1 => \N__4887\,
            in2 => \N__4875\,
            in3 => \N__4848\,
            lcout => \arse.g0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuresetoutreg_RNO_5_LC_24_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__4824\,
            in1 => \N__4811\,
            in2 => \N__4764\,
            in3 => \N__4736\,
            lcout => \arse.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.seven_LC_26_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4710\,
            lcout => \arse.divseven.sevenZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5391\,
            ce => \N__5352\,
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_2_LC_26_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110100000"
        )
    port map (
            in0 => \N__5437\,
            in1 => \N__5161\,
            in2 => \N__5196\,
            in3 => \N__5492\,
            lcout => \arse.divseven.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_0_LC_26_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010101010101"
        )
    port map (
            in0 => \N__5436\,
            in1 => \N__5157\,
            in2 => \N__5195\,
            in3 => \N__5491\,
            lcout => \arse.divseven.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.counter_1_LC_26_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001101001100"
        )
    port map (
            in0 => \N__5490\,
            in1 => \N__5187\,
            in2 => \N__5163\,
            in3 => \N__5438\,
            lcout => \arse.divseven.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.seven_RNO_LC_26_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__5489\,
            in1 => \N__5186\,
            in2 => \N__5162\,
            in3 => \N__5435\,
            lcout => \arse.divseven.N_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceup.out_e_0_LC_26_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5340\,
            lcout => debouncedup,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5308\,
            ce => \N__5241\,
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_RNO_0_0_LC_27_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__5434\,
            in1 => \N__5207\,
            in2 => \N__5194\,
            in3 => \N__5487\,
            lcout => OPEN,
            ltout => \arse.divseven.dout_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_0_LC_27_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__5488\,
            in1 => \_gnd_net_\,
            in2 => \N__5220\,
            in3 => \N__5152\,
            lcout => \arse.divseven.doutZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.divseven.dout_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_RNO_0_1_LC_27_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5185\,
            in2 => \_gnd_net_\,
            in3 => \N__5153\,
            lcout => \arse.divseven.un1_dout_2_sqmuxa_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounceconsolereset.out_RNI1B6C_LC_29_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5548\,
            lcout => debouncedconsolereset_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.cpuclkreset_LC_30_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__5698\,
            in1 => \N__5614\,
            in2 => \_gnd_net_\,
            in3 => \N__5133\,
            lcout => \arse.cpuclkresetZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.cpuclkresetC_net\,
            ce => 'H',
            sr => \N__5122\
        );

    \arse.diveight.counter_2_LC_31_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__5671\,
            in1 => \N__5607\,
            in2 => \N__5648\,
            in3 => \N__5579\,
            lcout => \arse.diveight.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_0_LC_31_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5667\,
            in2 => \_gnd_net_\,
            in3 => \N__5605\,
            lcout => \arse.diveight.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.counter_1_LC_31_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__5606\,
            in1 => \_gnd_net_\,
            in2 => \N__5673\,
            in3 => \N__5641\,
            lcout => \arse.diveight.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.apusynclatched_LC_32_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__5742\,
            in1 => \N__5684\,
            in2 => \_gnd_net_\,
            in3 => \N__5556\,
            lcout => \arse.apusynclatchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.apusynclatchedC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_1_LC_32_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__5672\,
            in1 => \N__5621\,
            in2 => \N__5649\,
            in3 => \N__5580\,
            lcout => \arse.diveight.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.diveight.dout_0_LC_32_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5622\,
            in2 => \_gnd_net_\,
            in3 => \N__5578\,
            lcout => \arse.diveight.doutZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.diveight.dout_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.apuresetoutreg_LC_32_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5555\,
            lcout => \arse.apuresetoutregZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVarse.diveight.dout_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \arse.divseven.dout_1_LC_32_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011110011001100"
        )
    port map (
            in0 => \N__5412\,
            in1 => \N__5502\,
            in2 => \N__5463\,
            in3 => \N__5445\,
            lcout => \arse.divseven.doutZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5394\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
