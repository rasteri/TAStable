// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 21 2024 23:56:49

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    masterreset,
    led4,
    lcol3,
    led5,
    lcol2,
    led6,
    led2,
    lcol1,
    deldn,
    cpuclk,
    apureset,
    altreset,
    led7,
    led3,
    lcol4,
    delup,
    cpureset,
    apusync,
    PACKAGEPIN,
    led8,
    led1,
    consolereset,
    apuclk);

    input masterreset;
    output led4;
    output lcol3;
    output led5;
    output lcol2;
    output led6;
    output led2;
    output lcol1;
    input deldn;
    output cpuclk;
    output apureset;
    input altreset;
    output led7;
    output led3;
    output lcol4;
    input delup;
    output cpureset;
    input apusync;
    input PACKAGEPIN;
    output led8;
    output led1;
    input consolereset;
    output apuclk;

    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6019;
    wire N__6018;
    wire N__6017;
    wire N__6010;
    wire N__6009;
    wire N__6008;
    wire N__6001;
    wire N__6000;
    wire N__5999;
    wire N__5992;
    wire N__5991;
    wire N__5990;
    wire N__5983;
    wire N__5982;
    wire N__5981;
    wire N__5974;
    wire N__5973;
    wire N__5972;
    wire N__5965;
    wire N__5964;
    wire N__5963;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5947;
    wire N__5946;
    wire N__5945;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5929;
    wire N__5928;
    wire N__5927;
    wire N__5920;
    wire N__5919;
    wire N__5918;
    wire N__5911;
    wire N__5910;
    wire N__5909;
    wire N__5902;
    wire N__5901;
    wire N__5900;
    wire N__5893;
    wire N__5892;
    wire N__5891;
    wire N__5884;
    wire N__5883;
    wire N__5882;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5866;
    wire N__5865;
    wire N__5864;
    wire N__5857;
    wire N__5856;
    wire N__5855;
    wire N__5848;
    wire N__5847;
    wire N__5846;
    wire N__5839;
    wire N__5838;
    wire N__5837;
    wire N__5830;
    wire N__5829;
    wire N__5828;
    wire N__5811;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5768;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5751;
    wire N__5750;
    wire N__5749;
    wire N__5748;
    wire N__5747;
    wire N__5746;
    wire N__5745;
    wire N__5744;
    wire N__5743;
    wire N__5742;
    wire N__5741;
    wire N__5740;
    wire N__5739;
    wire N__5738;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5690;
    wire N__5689;
    wire N__5688;
    wire N__5685;
    wire N__5684;
    wire N__5683;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5616;
    wire N__5615;
    wire N__5614;
    wire N__5613;
    wire N__5612;
    wire N__5611;
    wire N__5610;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5594;
    wire N__5589;
    wire N__5588;
    wire N__5587;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5575;
    wire N__5572;
    wire N__5571;
    wire N__5566;
    wire N__5563;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5529;
    wire N__5520;
    wire N__5517;
    wire N__5516;
    wire N__5515;
    wire N__5514;
    wire N__5513;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5496;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5470;
    wire N__5469;
    wire N__5464;
    wire N__5459;
    wire N__5454;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5413;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5388;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5369;
    wire N__5368;
    wire N__5365;
    wire N__5360;
    wire N__5355;
    wire N__5354;
    wire N__5353;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5341;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5315;
    wire N__5314;
    wire N__5313;
    wire N__5312;
    wire N__5311;
    wire N__5308;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5283;
    wire N__5282;
    wire N__5279;
    wire N__5274;
    wire N__5271;
    wire N__5264;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5240;
    wire N__5239;
    wire N__5238;
    wire N__5235;
    wire N__5228;
    wire N__5225;
    wire N__5220;
    wire N__5217;
    wire N__5208;
    wire N__5207;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5171;
    wire N__5170;
    wire N__5167;
    wire N__5162;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5144;
    wire N__5139;
    wire N__5138;
    wire N__5135;
    wire N__5134;
    wire N__5131;
    wire N__5126;
    wire N__5121;
    wire N__5120;
    wire N__5119;
    wire N__5116;
    wire N__5111;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5067;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5055;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5043;
    wire N__5042;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5027;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__4998;
    wire N__4997;
    wire N__4996;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4838;
    wire N__4835;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4802;
    wire N__4797;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4751;
    wire N__4750;
    wire N__4749;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4726;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4710;
    wire N__4707;
    wire N__4706;
    wire N__4703;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4695;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4677;
    wire N__4674;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4603;
    wire N__4602;
    wire N__4601;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4597;
    wire N__4596;
    wire N__4595;
    wire N__4594;
    wire N__4593;
    wire N__4592;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4541;
    wire N__4540;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4518;
    wire N__4515;
    wire N__4514;
    wire N__4513;
    wire N__4512;
    wire N__4511;
    wire N__4510;
    wire N__4509;
    wire N__4508;
    wire N__4507;
    wire N__4506;
    wire N__4505;
    wire N__4504;
    wire N__4503;
    wire N__4502;
    wire N__4501;
    wire N__4500;
    wire N__4499;
    wire N__4498;
    wire N__4497;
    wire N__4496;
    wire N__4495;
    wire N__4494;
    wire N__4493;
    wire N__4492;
    wire N__4491;
    wire N__4490;
    wire N__4489;
    wire N__4488;
    wire N__4487;
    wire N__4484;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4415;
    wire N__4414;
    wire N__4413;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4405;
    wire N__4404;
    wire N__4403;
    wire N__4400;
    wire N__4395;
    wire N__4390;
    wire N__4385;
    wire N__4384;
    wire N__4381;
    wire N__4376;
    wire N__4375;
    wire N__4374;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4326;
    wire N__4323;
    wire N__4322;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4304;
    wire N__4303;
    wire N__4300;
    wire N__4299;
    wire N__4296;
    wire N__4295;
    wire N__4294;
    wire N__4289;
    wire N__4286;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4260;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4239;
    wire N__4236;
    wire N__4231;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4206;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4190;
    wire N__4187;
    wire N__4186;
    wire N__4185;
    wire N__4182;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4118;
    wire N__4115;
    wire N__4114;
    wire N__4111;
    wire N__4110;
    wire N__4109;
    wire N__4106;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4090;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4053;
    wire N__4052;
    wire N__4051;
    wire N__4050;
    wire N__4049;
    wire N__4048;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4019;
    wire N__4018;
    wire N__4015;
    wire N__4010;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3980;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3965;
    wire N__3960;
    wire N__3957;
    wire N__3956;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3933;
    wire N__3932;
    wire N__3931;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3903;
    wire N__3902;
    wire N__3899;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3882;
    wire N__3879;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3836;
    wire N__3833;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3819;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3745;
    wire N__3740;
    wire N__3739;
    wire N__3738;
    wire N__3737;
    wire N__3736;
    wire N__3733;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3725;
    wire N__3722;
    wire N__3721;
    wire N__3720;
    wire N__3719;
    wire N__3716;
    wire N__3711;
    wire N__3710;
    wire N__3709;
    wire N__3706;
    wire N__3701;
    wire N__3698;
    wire N__3693;
    wire N__3692;
    wire N__3691;
    wire N__3688;
    wire N__3687;
    wire N__3686;
    wire N__3683;
    wire N__3678;
    wire N__3673;
    wire N__3672;
    wire N__3667;
    wire N__3666;
    wire N__3661;
    wire N__3660;
    wire N__3659;
    wire N__3658;
    wire N__3657;
    wire N__3654;
    wire N__3645;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3621;
    wire N__3616;
    wire N__3613;
    wire N__3608;
    wire N__3591;
    wire N__3588;
    wire N__3587;
    wire N__3586;
    wire N__3583;
    wire N__3582;
    wire N__3581;
    wire N__3580;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3572;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3561;
    wire N__3560;
    wire N__3559;
    wire N__3558;
    wire N__3557;
    wire N__3556;
    wire N__3555;
    wire N__3554;
    wire N__3553;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3517;
    wire N__3514;
    wire N__3509;
    wire N__3508;
    wire N__3505;
    wire N__3500;
    wire N__3497;
    wire N__3492;
    wire N__3489;
    wire N__3488;
    wire N__3479;
    wire N__3478;
    wire N__3477;
    wire N__3476;
    wire N__3475;
    wire N__3474;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3458;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3437;
    wire N__3432;
    wire N__3427;
    wire N__3420;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3366;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3347;
    wire N__3344;
    wire N__3343;
    wire N__3342;
    wire N__3339;
    wire N__3336;
    wire N__3331;
    wire N__3328;
    wire N__3321;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3313;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3213;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3201;
    wire N__3200;
    wire N__3197;
    wire N__3196;
    wire N__3193;
    wire N__3188;
    wire N__3183;
    wire N__3182;
    wire N__3181;
    wire N__3180;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3162;
    wire N__3161;
    wire N__3158;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3141;
    wire N__3138;
    wire N__3137;
    wire N__3136;
    wire N__3135;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3117;
    wire N__3114;
    wire N__3113;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3096;
    wire N__3095;
    wire N__3092;
    wire N__3091;
    wire N__3088;
    wire N__3087;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2987;
    wire N__2986;
    wire N__2983;
    wire N__2978;
    wire N__2977;
    wire N__2976;
    wire N__2975;
    wire N__2974;
    wire N__2973;
    wire N__2972;
    wire N__2971;
    wire N__2970;
    wire N__2969;
    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2965;
    wire N__2964;
    wire N__2963;
    wire N__2958;
    wire N__2951;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2929;
    wire N__2922;
    wire N__2919;
    wire N__2904;
    wire N__2903;
    wire N__2900;
    wire N__2899;
    wire N__2896;
    wire N__2895;
    wire N__2894;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2877;
    wire N__2874;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2682;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2670;
    wire N__2667;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2655;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2643;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2631;
    wire N__2628;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2591;
    wire N__2590;
    wire N__2587;
    wire N__2582;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2563;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2541;
    wire N__2538;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2526;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2502;
    wire N__2501;
    wire N__2500;
    wire N__2499;
    wire N__2492;
    wire N__2489;
    wire N__2486;
    wire N__2481;
    wire N__2480;
    wire N__2479;
    wire N__2476;
    wire N__2471;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2457;
    wire N__2454;
    wire N__2451;
    wire N__2448;
    wire N__2445;
    wire N__2442;
    wire N__2441;
    wire N__2438;
    wire N__2435;
    wire N__2430;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2418;
    wire N__2415;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2400;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2388;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2376;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2364;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2352;
    wire N__2349;
    wire N__2346;
    wire N__2343;
    wire N__2340;
    wire N__2337;
    wire N__2334;
    wire N__2331;
    wire N__2328;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2316;
    wire N__2313;
    wire N__2310;
    wire N__2307;
    wire N__2304;
    wire N__2301;
    wire N__2298;
    wire N__2295;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2274;
    wire N__2271;
    wire N__2268;
    wire N__2265;
    wire N__2262;
    wire N__2259;
    wire N__2256;
    wire N__2253;
    wire N__2250;
    wire N__2247;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2211;
    wire N__2208;
    wire N__2205;
    wire N__2202;
    wire N__2199;
    wire N__2196;
    wire \arse.un1_io_0_1_g ;
    wire \top_pll_nrtthrth.PLLOUTCORE ;
    wire GNDG0;
    wire \arse.divseven.io_0_D_IN_0 ;
    wire VCCG0;
    wire masterreset_c_i;
    wire bfn_15_18_0_;
    wire \debounceup.un3_counter_1_cry_1 ;
    wire \debounceup.un3_counter_1_cry_2 ;
    wire \debounceup.un3_counter_1_cry_3 ;
    wire bfn_15_23_0_;
    wire \arses.un2_counter_cry_1 ;
    wire \arses.un2_counter_cry_2 ;
    wire \arses.un2_counter_cry_3 ;
    wire \arses.un2_counter_cry_4 ;
    wire \arses.un2_counter_cry_5 ;
    wire \arses.un2_counter_cry_6 ;
    wire \arses.un2_counter_cry_7 ;
    wire \arses.un2_counter_cry_8 ;
    wire bfn_15_24_0_;
    wire \arses.un2_counter_cry_9 ;
    wire \arses.un2_counter_cry_10 ;
    wire \arses.un2_counter_cry_11 ;
    wire \arses.un2_counter_cry_12 ;
    wire \arses.un2_counter_cry_13 ;
    wire lcol4_c;
    wire GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO;
    wire \debounceup.counterZ0Z_3 ;
    wire \debounceup.counter19_2_cascade_ ;
    wire \debounceup.counter_RNO_0_0_2 ;
    wire \debounceup.counter19_cascade_ ;
    wire \debounceup.counterZ0Z_2 ;
    wire \debounceup.counterZ0Z_4 ;
    wire \debounceup.counter19_2 ;
    wire \dig2.m18_bm_cascade_ ;
    wire leds_1_i_1;
    wire \arses.counterZ0Z_7 ;
    wire \arses.counterZ0Z_6 ;
    wire \arses.counterZ0Z_5 ;
    wire \arses.counterZ0Z_8 ;
    wire \arses.counterZ0Z_3 ;
    wire \arses.counterZ0Z_2 ;
    wire \arses.counterZ0Z_4 ;
    wire \arses.un1_counterlto4_2_cascade_ ;
    wire \arses.un1_counterlto8_2 ;
    wire \arses.counterZ0Z_11 ;
    wire \arses.counterZ0Z_10 ;
    wire \arses.un1_counterlt11_cascade_ ;
    wire \arses.counterZ0Z_9 ;
    wire \arses.counterZ0Z_14 ;
    wire \arses.counterZ0Z_13 ;
    wire \arses.un1_counterlt13_0_cascade_ ;
    wire \arses.counterZ0Z_12 ;
    wire arses_counter8_cascade_;
    wire \arses.clock_out_RNIR6ERZ0Z_0 ;
    wire \arses.counterZ0Z_1 ;
    wire \arses.counterZ0Z_0 ;
    wire lcol3_c;
    wire \dig2.m13_am_cascade_ ;
    wire \dig2.leds_17_i_0_ns_1_1 ;
    wire \dig2.m18_am ;
    wire leds_1_i_3;
    wire \dig2.m13_bm ;
    wire \dig2.N_42 ;
    wire \dig2.m69_am ;
    wire \dig2.m69_bm ;
    wire leds_1_i_0_2;
    wire \dig2.N_78 ;
    wire \dig2.N_76 ;
    wire leds_1_i_0_3;
    wire \dig2.m39_ns_1_cascade_ ;
    wire \dig2.N_40 ;
    wire \dig2.i3_mux ;
    wire \dig2.N_59 ;
    wire \dig2.leds_17_i_ns_1_2 ;
    wire consolereset_c;
    wire altreset_c;
    wire \debounceconsolereset.out_RNOZ0Z_0_cascade_ ;
    wire clock_out_RNIR6ER;
    wire clock_out_RNIR6ER_cascade_;
    wire arses_counter8;
    wire slowclk;
    wire \dig2.m54_am ;
    wire leds_1_i_0_1;
    wire \dig2.m75_ns_1 ;
    wire bfn_20_17_0_;
    wire \debounceconsolereset.counter_RNO_0Z0Z_2 ;
    wire \debounceconsolereset.un3_counter_1_cry_1 ;
    wire \debounceconsolereset.un3_counter_1_cry_2 ;
    wire \debounceconsolereset.un3_counter_1_cry_3 ;
    wire \debounceconsolereset.counterZ0Z_3 ;
    wire \debounceconsolereset.counterZ0Z_2 ;
    wire \debounceconsolereset.counter19_2 ;
    wire \debounceconsolereset.counterZ0Z_4 ;
    wire \debounceconsolereset.counterZ0Z_1 ;
    wire \debounceconsolereset.counter19_2_cascade_ ;
    wire \debounceconsolereset.counterZ0Z_0 ;
    wire \debounceconsolereset.counter19 ;
    wire col_1_1;
    wire \dig2.m54_bm ;
    wire \dig2.leds_17_i_ns_1_1 ;
    wire \debounceup.counterZ0Z_0 ;
    wire \debounceup.counterZ0Z_1 ;
    wire \dig2.m49_bm ;
    wire \dig2.m49_am ;
    wire \dig2.m33_am ;
    wire \dig2.m33_bm_cascade_ ;
    wire leds_1_i_2;
    wire \dig2.N_25_cascade_ ;
    wire \dig2.leds_17_i_0_ns_1_2 ;
    wire \dig2.i2_mux ;
    wire lcol1_c;
    wire colZ0Z_1;
    wire colZ0Z_0;
    wire lcol2_c;
    wire \debouncedn.counter19_2_cascade_ ;
    wire \debouncedn.counter19_cascade_ ;
    wire bfn_24_17_0_;
    wire \debouncedn.counterZ0Z_2 ;
    wire \debouncedn.counter_RNO_0_1_2 ;
    wire \debouncedn.un3_counter_1_cry_1 ;
    wire \debouncedn.counterZ0Z_3 ;
    wire \debouncedn.un3_counter_1_cry_2 ;
    wire \debouncedn.counter19_2 ;
    wire \debouncedn.un3_counter_1_cry_3 ;
    wire \debouncedn.counterZ0Z_4 ;
    wire \debouncedn.counterZ0Z_0 ;
    wire \debouncedn.counterZ0Z_1 ;
    wire \debouncedn.counter19 ;
    wire deldn_c;
    wire CONSTANT_ONE_NET;
    wire bfn_27_10_0_;
    wire un1_delayConstant_cry_0;
    wire un1_delayConstant_cry_1;
    wire un1_delayConstant_cry_2;
    wire delayConstantZ0Z_4;
    wire un1_delayConstant_cry_3;
    wire delayConstantZ0Z_5;
    wire un1_delayConstant_cry_4;
    wire delayConstantZ0Z_6;
    wire un1_delayConstant_cry_5;
    wire un1_delayConstant_cry_6;
    wire delayConstantZ0Z_7;
    wire masterreset_c_i_g;
    wire olddnZ0;
    wire debounceddn;
    wire olddn_RNIEENHZ0_cascade_;
    wire olddn_RNIM5BH1Z0Z_0;
    wire olddn_RNIM5BH1Z0Z_3;
    wire olddn_RNIM5BH1Z0Z_1;
    wire masterreset_c;
    wire delayConstant17_i_cascade_;
    wire un1_delayConstant_cry_0_c_RNOZ0;
    wire olddn_RNIM5BH1Z0Z_4;
    wire olddn_RNIM5BHZ0Z1;
    wire olddn_RNIEENHZ0;
    wire delayConstant17_i;
    wire olddn_RNIM5BH1Z0Z_2;
    wire oldupZ0;
    wire \debounceup.counter19 ;
    wire delup_c;
    wire N_111_g;
    wire debouncedup;
    wire PACKAGEPIN_0_c_g;
    wire bfn_29_7_0_;
    wire \arse.un1_cpuresetcount_1_cry_0 ;
    wire \arse.un1_cpuresetcount_1_cry_1 ;
    wire \arse.un1_cpuresetcount_1_cry_2 ;
    wire \arse.un1_cpuresetcount_1_cry_3 ;
    wire \arse.un1_cpuresetcount_1_cry_4 ;
    wire \arse.un1_cpuresetcount_1_cry_5 ;
    wire \arse.un1_cpuresetcount_1_cry_6 ;
    wire \INVarse.cpuresetcount_0C_net ;
    wire \arse.cpuresetoutregZ0 ;
    wire \INVarse.cpuresetoutregC_net ;
    wire \arse.m8_2_cascade_ ;
    wire \arse.cpuresetcountZ0Z_0 ;
    wire \arse.cpuresetcountZ0Z_5 ;
    wire \arse.cpuresetcountZ0Z_1 ;
    wire \arse.cpuresetcountZ0Z_2 ;
    wire \arse.m12_2_cascade_ ;
    wire \arse.cpuresetcountZ0Z_4 ;
    wire \arse.cpuresetoutreg_1_sqmuxa ;
    wire \arse.cpuresetcountZ0Z_7 ;
    wire \arse.cpuresetcountZ0Z_6 ;
    wire \arse.cpuresetcountZ0Z_3 ;
    wire \arse.m4_e_2 ;
    wire \arse.cpuclkreset_1_sqmuxa ;
    wire \INVarse.cpuclkresetC_net ;
    wire debouncedconsolereset_i;
    wire \INVarse.diveight.dout_0C_net ;
    wire delayConstantZ0Z_3;
    wire arse_diveight_N_123_0_cascade_;
    wire delayConstantZ0Z_2;
    wire delayConstantZ0Z_1;
    wire arse_cpuclkreset;
    wire apusync_c;
    wire \arse.apusynclatchedZ0 ;
    wire \INVarse.apusynclatchedC_net ;
    wire \arse.diveight.doutZ0Z_0 ;
    wire \arse.diveight.dout_i_0 ;
    wire \arse.diveight.dout_i_1 ;
    wire debouncedconsolereset;
    wire \arse.apuresetoutregZ0 ;
    wire \INVarse.apuresetoutregC_net ;
    wire arse_diveight_counter_1;
    wire arse_diveight_counter_0;
    wire delayConstantZ0Z_0;
    wire arse_diveight_counter_2;
    wire \arse.diveight.doutZ0Z_1 ;
    wire \arse.diveight.cpuclkreset_i ;
    wire \arse.divseven.counterZ0Z_1 ;
    wire \arse.divseven.counterZ0Z_0 ;
    wire \INVarse.divseven.dout_0C_net ;
    wire \arse.divseven.doutZ0Z_0 ;
    wire \arse.divseven.dout_i_0 ;
    wire \arse.divseven.counterZ0Z_2 ;
    wire PLLOUTCORE_g;
    wire \arse.divseven.doutZ0Z_1 ;
    wire \arse.divseven.dout_i_1 ;
    wire _gnd_net_;

    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .TEST_MODE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FILTER_RANGE=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_RELATIVE=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVR=4'b0000;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVQ=3'b010;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DIVF=7'b0011111;
    defparam \top_pll_nrtthrth.top_pll_nrtthrth_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \top_pll_nrtthrth.top_pll_nrtthrth_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\top_pll_nrtthrth.PLLOUTCORE ),
            .REFERENCECLK(N__2304),
            .RESETB(N__4878),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF PACKAGEPIN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6028),
            .GLOBALBUFFEROUTPUT(PACKAGEPIN_0_c_g));
    IO_PAD PACKAGEPIN_ibuf_gb_io_iopad (
            .OE(N__6030),
            .DIN(N__6029),
            .DOUT(N__6028),
            .PACKAGEPIN(PACKAGEPIN));
    defparam PACKAGEPIN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam PACKAGEPIN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO PACKAGEPIN_ibuf_gb_io_preio (
            .PADOEN(N__6030),
            .PADOUT(N__6029),
            .PADIN(N__6028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD masterreset_ibuf_iopad (
            .OE(N__6019),
            .DIN(N__6018),
            .DOUT(N__6017),
            .PACKAGEPIN(masterreset));
    defparam masterreset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam masterreset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO masterreset_ibuf_preio (
            .PADOEN(N__6019),
            .PADOUT(N__6018),
            .PADIN(N__6017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(masterreset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led3_obuf_iopad (
            .OE(N__6010),
            .DIN(N__6009),
            .DOUT(N__6008),
            .PACKAGEPIN(led3));
    defparam led3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led3_obuf_preio (
            .PADOEN(N__6010),
            .PADOUT(N__6009),
            .PADIN(N__6008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2820),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.divseven.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.divseven.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.divseven.io_0_iopad  (
            .OE(N__6001),
            .DIN(N__6000),
            .DOUT(N__5999),
            .PACKAGEPIN(apuclk));
    defparam \arse.divseven.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.divseven.io_0_preio  (
            .PADOEN(N__6001),
            .PADOUT(N__6000),
            .PADIN(N__5999),
            .CLOCKENABLE(),
            .DOUT1(N__5697),
            .OUTPUTENABLE(N__3832),
            .DIN0(\arse.divseven.io_0_D_IN_0 ),
            .DOUT0(N__5778),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5738));
    defparam \arse.io_1_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.io_1_iopad .PULLUP=1'b0;
    IO_PAD \arse.io_1_iopad  (
            .OE(N__5992),
            .DIN(N__5991),
            .DOUT(N__5990),
            .PACKAGEPIN(cpureset));
    defparam \arse.io_1_preio .PIN_TYPE=6'b010101;
    PRE_IO \arse.io_1_preio  (
            .PADOEN(N__5992),
            .PADOUT(N__5991),
            .PADIN(N__5990),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4896),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5748));
    IO_PAD lcol3_obuf_iopad (
            .OE(N__5983),
            .DIN(N__5982),
            .DOUT(N__5981),
            .PACKAGEPIN(lcol3));
    defparam lcol3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol3_obuf_preio (
            .PADOEN(N__5983),
            .PADOUT(N__5982),
            .PADIN(N__5981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2556),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD deldn_ibuf_iopad (
            .OE(N__5974),
            .DIN(N__5973),
            .DOUT(N__5972),
            .PACKAGEPIN(deldn));
    defparam deldn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam deldn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO deldn_ibuf_preio (
            .PADOEN(N__5974),
            .PADOUT(N__5973),
            .PADIN(N__5972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(deldn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led2_obuf_iopad (
            .OE(N__5965),
            .DIN(N__5964),
            .DOUT(N__5963),
            .PACKAGEPIN(led2));
    defparam led2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led2_obuf_preio (
            .PADOEN(N__5965),
            .PADOUT(N__5964),
            .PADIN(N__5963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delup_ibuf_iopad (
            .OE(N__5956),
            .DIN(N__5955),
            .DOUT(N__5954),
            .PACKAGEPIN(delup));
    defparam delup_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delup_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delup_ibuf_preio (
            .PADOEN(N__5956),
            .PADOUT(N__5955),
            .PADIN(N__5954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delup_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led6_obuf_iopad (
            .OE(N__5947),
            .DIN(N__5946),
            .DOUT(N__5945),
            .PACKAGEPIN(led6));
    defparam led6_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led6_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led6_obuf_preio (
            .PADOEN(N__5947),
            .PADOUT(N__5946),
            .PADIN(N__5945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led8_obuf_iopad (
            .OE(N__5938),
            .DIN(N__5937),
            .DOUT(N__5936),
            .PACKAGEPIN(led8));
    defparam led8_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led8_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led8_obuf_preio (
            .PADOEN(N__5938),
            .PADOUT(N__5937),
            .PADIN(N__5936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD altreset_ibuf_iopad (
            .OE(N__5929),
            .DIN(N__5928),
            .DOUT(N__5927),
            .PACKAGEPIN(altreset));
    defparam altreset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam altreset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO altreset_ibuf_preio (
            .PADOEN(N__5929),
            .PADOUT(N__5928),
            .PADIN(N__5927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(altreset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led4_obuf_iopad (
            .OE(N__5920),
            .DIN(N__5919),
            .DOUT(N__5918),
            .PACKAGEPIN(led4));
    defparam led4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led4_obuf_preio (
            .PADOEN(N__5920),
            .PADOUT(N__5919),
            .PADIN(N__5918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2784),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.io_0_iopad  (
            .OE(N__5911),
            .DIN(N__5910),
            .DOUT(N__5909),
            .PACKAGEPIN(apureset));
    defparam \arse.io_0_preio .PIN_TYPE=6'b010101;
    PRE_IO \arse.io_0_preio  (
            .PADOEN(N__5911),
            .PADOUT(N__5910),
            .PADIN(N__5909),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5376),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5744));
    IO_PAD lcol4_obuf_iopad (
            .OE(N__5902),
            .DIN(N__5901),
            .DOUT(N__5900),
            .PACKAGEPIN(lcol4));
    defparam lcol4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol4_obuf_preio (
            .PADOEN(N__5902),
            .PADOUT(N__5901),
            .PADIN(N__5900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2322),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam \arse.diveight.io_0_iopad .IO_STANDARD="SB_LVCMOS";
    defparam \arse.diveight.io_0_iopad .PULLUP=1'b0;
    IO_PAD \arse.diveight.io_0_iopad  (
            .OE(N__5893),
            .DIN(N__5892),
            .DOUT(N__5891),
            .PACKAGEPIN(cpuclk));
    defparam \arse.diveight.io_0_preio .PIN_TYPE=6'b100001;
    PRE_IO \arse.diveight.io_0_preio  (
            .PADOEN(N__5893),
            .PADOUT(N__5892),
            .PADIN(N__5891),
            .CLOCKENABLE(),
            .DOUT1(N__5430),
            .OUTPUTENABLE(N__3840),
            .DIN0(),
            .DOUT0(N__5436),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK(N__5744));
    IO_PAD led5_obuf_iopad (
            .OE(N__5884),
            .DIN(N__5883),
            .DOUT(N__5882),
            .PACKAGEPIN(led5));
    defparam led5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led5_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led5_obuf_preio (
            .PADOEN(N__5884),
            .PADOUT(N__5883),
            .PADIN(N__5882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3836),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD consolereset_ibuf_iopad (
            .OE(N__5875),
            .DIN(N__5874),
            .DOUT(N__5873),
            .PACKAGEPIN(consolereset));
    defparam consolereset_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam consolereset_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO consolereset_ibuf_preio (
            .PADOEN(N__5875),
            .PADOUT(N__5874),
            .PADIN(N__5873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(consolereset_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol2_obuf_iopad (
            .OE(N__5866),
            .DIN(N__5865),
            .DOUT(N__5864),
            .PACKAGEPIN(lcol2));
    defparam lcol2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol2_obuf_preio (
            .PADOEN(N__5866),
            .PADOUT(N__5865),
            .PADIN(N__5864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3405),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led1_obuf_iopad (
            .OE(N__5857),
            .DIN(N__5856),
            .DOUT(N__5855),
            .PACKAGEPIN(led1));
    defparam led1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led1_obuf_preio (
            .PADOEN(N__5857),
            .PADOUT(N__5856),
            .PADIN(N__5855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3819),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD apusync_ibuf_iopad (
            .OE(N__5848),
            .DIN(N__5847),
            .DOUT(N__5846),
            .PACKAGEPIN(apusync));
    defparam apusync_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam apusync_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO apusync_ibuf_preio (
            .PADOEN(N__5848),
            .PADOUT(N__5847),
            .PADIN(N__5846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(apusync_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led7_obuf_iopad (
            .OE(N__5839),
            .DIN(N__5838),
            .DOUT(N__5837),
            .PACKAGEPIN(led7));
    defparam led7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam led7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO led7_obuf_preio (
            .PADOEN(N__5839),
            .PADOUT(N__5838),
            .PADIN(N__5837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3273),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD lcol1_obuf_iopad (
            .OE(N__5830),
            .DIN(N__5829),
            .DOUT(N__5828),
            .PACKAGEPIN(lcol1));
    defparam lcol1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam lcol1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO lcol1_obuf_preio (
            .PADOEN(N__5830),
            .PADOUT(N__5829),
            .PADIN(N__5828),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3768),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1401 (
            .O(N__5811),
            .I(N__5807));
    InMux I__1400 (
            .O(N__5810),
            .I(N__5804));
    LocalMux I__1399 (
            .O(N__5807),
            .I(\arse.divseven.counterZ0Z_1 ));
    LocalMux I__1398 (
            .O(N__5804),
            .I(\arse.divseven.counterZ0Z_1 ));
    InMux I__1397 (
            .O(N__5799),
            .I(N__5790));
    InMux I__1396 (
            .O(N__5798),
            .I(N__5790));
    InMux I__1395 (
            .O(N__5797),
            .I(N__5790));
    LocalMux I__1394 (
            .O(N__5790),
            .I(\arse.divseven.counterZ0Z_0 ));
    CascadeMux I__1393 (
            .O(N__5787),
            .I(N__5784));
    InMux I__1392 (
            .O(N__5784),
            .I(N__5781));
    LocalMux I__1391 (
            .O(N__5781),
            .I(\arse.divseven.doutZ0Z_0 ));
    IoInMux I__1390 (
            .O(N__5778),
            .I(N__5775));
    LocalMux I__1389 (
            .O(N__5775),
            .I(\arse.divseven.dout_i_0 ));
    InMux I__1388 (
            .O(N__5772),
            .I(N__5769));
    LocalMux I__1387 (
            .O(N__5769),
            .I(N__5764));
    InMux I__1386 (
            .O(N__5768),
            .I(N__5761));
    InMux I__1385 (
            .O(N__5767),
            .I(N__5758));
    Odrv12 I__1384 (
            .O(N__5764),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__1383 (
            .O(N__5761),
            .I(\arse.divseven.counterZ0Z_2 ));
    LocalMux I__1382 (
            .O(N__5758),
            .I(\arse.divseven.counterZ0Z_2 ));
    ClkMux I__1381 (
            .O(N__5751),
            .I(N__5709));
    ClkMux I__1380 (
            .O(N__5750),
            .I(N__5709));
    ClkMux I__1379 (
            .O(N__5749),
            .I(N__5709));
    ClkMux I__1378 (
            .O(N__5748),
            .I(N__5709));
    ClkMux I__1377 (
            .O(N__5747),
            .I(N__5709));
    ClkMux I__1376 (
            .O(N__5746),
            .I(N__5709));
    ClkMux I__1375 (
            .O(N__5745),
            .I(N__5709));
    ClkMux I__1374 (
            .O(N__5744),
            .I(N__5709));
    ClkMux I__1373 (
            .O(N__5743),
            .I(N__5709));
    ClkMux I__1372 (
            .O(N__5742),
            .I(N__5709));
    ClkMux I__1371 (
            .O(N__5741),
            .I(N__5709));
    ClkMux I__1370 (
            .O(N__5740),
            .I(N__5709));
    ClkMux I__1369 (
            .O(N__5739),
            .I(N__5709));
    ClkMux I__1368 (
            .O(N__5738),
            .I(N__5709));
    GlobalMux I__1367 (
            .O(N__5709),
            .I(N__5706));
    gio2CtrlBuf I__1366 (
            .O(N__5706),
            .I(PLLOUTCORE_g));
    InMux I__1365 (
            .O(N__5703),
            .I(N__5700));
    LocalMux I__1364 (
            .O(N__5700),
            .I(\arse.divseven.doutZ0Z_1 ));
    IoInMux I__1363 (
            .O(N__5697),
            .I(N__5694));
    LocalMux I__1362 (
            .O(N__5694),
            .I(\arse.divseven.dout_i_1 ));
    CascadeMux I__1361 (
            .O(N__5691),
            .I(N__5685));
    InMux I__1360 (
            .O(N__5690),
            .I(N__5678));
    InMux I__1359 (
            .O(N__5689),
            .I(N__5678));
    InMux I__1358 (
            .O(N__5688),
            .I(N__5675));
    InMux I__1357 (
            .O(N__5685),
            .I(N__5672));
    CascadeMux I__1356 (
            .O(N__5684),
            .I(N__5669));
    CascadeMux I__1355 (
            .O(N__5683),
            .I(N__5666));
    LocalMux I__1354 (
            .O(N__5678),
            .I(N__5659));
    LocalMux I__1353 (
            .O(N__5675),
            .I(N__5659));
    LocalMux I__1352 (
            .O(N__5672),
            .I(N__5659));
    InMux I__1351 (
            .O(N__5669),
            .I(N__5656));
    InMux I__1350 (
            .O(N__5666),
            .I(N__5653));
    Span4Mux_v I__1349 (
            .O(N__5659),
            .I(N__5650));
    LocalMux I__1348 (
            .O(N__5656),
            .I(N__5646));
    LocalMux I__1347 (
            .O(N__5653),
            .I(N__5643));
    Span4Mux_h I__1346 (
            .O(N__5650),
            .I(N__5640));
    CascadeMux I__1345 (
            .O(N__5649),
            .I(N__5637));
    Span4Mux_v I__1344 (
            .O(N__5646),
            .I(N__5634));
    Span12Mux_v I__1343 (
            .O(N__5643),
            .I(N__5631));
    Span4Mux_v I__1342 (
            .O(N__5640),
            .I(N__5628));
    InMux I__1341 (
            .O(N__5637),
            .I(N__5625));
    Odrv4 I__1340 (
            .O(N__5634),
            .I(delayConstantZ0Z_2));
    Odrv12 I__1339 (
            .O(N__5631),
            .I(delayConstantZ0Z_2));
    Odrv4 I__1338 (
            .O(N__5628),
            .I(delayConstantZ0Z_2));
    LocalMux I__1337 (
            .O(N__5625),
            .I(delayConstantZ0Z_2));
    InMux I__1336 (
            .O(N__5616),
            .I(N__5606));
    InMux I__1335 (
            .O(N__5615),
            .I(N__5603));
    InMux I__1334 (
            .O(N__5614),
            .I(N__5594));
    InMux I__1333 (
            .O(N__5613),
            .I(N__5594));
    InMux I__1332 (
            .O(N__5612),
            .I(N__5594));
    InMux I__1331 (
            .O(N__5611),
            .I(N__5594));
    InMux I__1330 (
            .O(N__5610),
            .I(N__5589));
    InMux I__1329 (
            .O(N__5609),
            .I(N__5589));
    LocalMux I__1328 (
            .O(N__5606),
            .I(N__5583));
    LocalMux I__1327 (
            .O(N__5603),
            .I(N__5580));
    LocalMux I__1326 (
            .O(N__5594),
            .I(N__5575));
    LocalMux I__1325 (
            .O(N__5589),
            .I(N__5575));
    InMux I__1324 (
            .O(N__5588),
            .I(N__5572));
    InMux I__1323 (
            .O(N__5587),
            .I(N__5566));
    InMux I__1322 (
            .O(N__5586),
            .I(N__5566));
    Span4Mux_h I__1321 (
            .O(N__5583),
            .I(N__5563));
    Span4Mux_v I__1320 (
            .O(N__5580),
            .I(N__5558));
    Span4Mux_v I__1319 (
            .O(N__5575),
            .I(N__5558));
    LocalMux I__1318 (
            .O(N__5572),
            .I(N__5555));
    CascadeMux I__1317 (
            .O(N__5571),
            .I(N__5552));
    LocalMux I__1316 (
            .O(N__5566),
            .I(N__5549));
    Span4Mux_h I__1315 (
            .O(N__5563),
            .I(N__5546));
    Sp12to4 I__1314 (
            .O(N__5558),
            .I(N__5543));
    Span4Mux_v I__1313 (
            .O(N__5555),
            .I(N__5540));
    InMux I__1312 (
            .O(N__5552),
            .I(N__5537));
    Span12Mux_v I__1311 (
            .O(N__5549),
            .I(N__5534));
    Sp12to4 I__1310 (
            .O(N__5546),
            .I(N__5529));
    Span12Mux_h I__1309 (
            .O(N__5543),
            .I(N__5529));
    Odrv4 I__1308 (
            .O(N__5540),
            .I(delayConstantZ0Z_1));
    LocalMux I__1307 (
            .O(N__5537),
            .I(delayConstantZ0Z_1));
    Odrv12 I__1306 (
            .O(N__5534),
            .I(delayConstantZ0Z_1));
    Odrv12 I__1305 (
            .O(N__5529),
            .I(delayConstantZ0Z_1));
    InMux I__1304 (
            .O(N__5520),
            .I(N__5517));
    LocalMux I__1303 (
            .O(N__5517),
            .I(N__5509));
    InMux I__1302 (
            .O(N__5516),
            .I(N__5506));
    InMux I__1301 (
            .O(N__5515),
            .I(N__5503));
    InMux I__1300 (
            .O(N__5514),
            .I(N__5496));
    InMux I__1299 (
            .O(N__5513),
            .I(N__5496));
    InMux I__1298 (
            .O(N__5512),
            .I(N__5496));
    Odrv4 I__1297 (
            .O(N__5509),
            .I(arse_cpuclkreset));
    LocalMux I__1296 (
            .O(N__5506),
            .I(arse_cpuclkreset));
    LocalMux I__1295 (
            .O(N__5503),
            .I(arse_cpuclkreset));
    LocalMux I__1294 (
            .O(N__5496),
            .I(arse_cpuclkreset));
    InMux I__1293 (
            .O(N__5487),
            .I(N__5484));
    LocalMux I__1292 (
            .O(N__5484),
            .I(apusync_c));
    CascadeMux I__1291 (
            .O(N__5481),
            .I(N__5477));
    InMux I__1290 (
            .O(N__5480),
            .I(N__5474));
    InMux I__1289 (
            .O(N__5477),
            .I(N__5471));
    LocalMux I__1288 (
            .O(N__5474),
            .I(N__5464));
    LocalMux I__1287 (
            .O(N__5471),
            .I(N__5464));
    InMux I__1286 (
            .O(N__5470),
            .I(N__5459));
    InMux I__1285 (
            .O(N__5469),
            .I(N__5459));
    Span4Mux_h I__1284 (
            .O(N__5464),
            .I(N__5454));
    LocalMux I__1283 (
            .O(N__5459),
            .I(N__5454));
    Span4Mux_v I__1282 (
            .O(N__5454),
            .I(N__5450));
    InMux I__1281 (
            .O(N__5453),
            .I(N__5447));
    Odrv4 I__1280 (
            .O(N__5450),
            .I(\arse.apusynclatchedZ0 ));
    LocalMux I__1279 (
            .O(N__5447),
            .I(\arse.apusynclatchedZ0 ));
    InMux I__1278 (
            .O(N__5442),
            .I(N__5439));
    LocalMux I__1277 (
            .O(N__5439),
            .I(\arse.diveight.doutZ0Z_0 ));
    IoInMux I__1276 (
            .O(N__5436),
            .I(N__5433));
    LocalMux I__1275 (
            .O(N__5433),
            .I(\arse.diveight.dout_i_0 ));
    IoInMux I__1274 (
            .O(N__5430),
            .I(N__5427));
    LocalMux I__1273 (
            .O(N__5427),
            .I(\arse.diveight.dout_i_1 ));
    InMux I__1272 (
            .O(N__5424),
            .I(N__5421));
    LocalMux I__1271 (
            .O(N__5421),
            .I(N__5417));
    InMux I__1270 (
            .O(N__5420),
            .I(N__5414));
    Span4Mux_s0_h I__1269 (
            .O(N__5417),
            .I(N__5408));
    LocalMux I__1268 (
            .O(N__5414),
            .I(N__5408));
    InMux I__1267 (
            .O(N__5413),
            .I(N__5405));
    Span4Mux_v I__1266 (
            .O(N__5408),
            .I(N__5402));
    LocalMux I__1265 (
            .O(N__5405),
            .I(N__5399));
    Span4Mux_v I__1264 (
            .O(N__5402),
            .I(N__5396));
    Span4Mux_v I__1263 (
            .O(N__5399),
            .I(N__5393));
    Sp12to4 I__1262 (
            .O(N__5396),
            .I(N__5388));
    Sp12to4 I__1261 (
            .O(N__5393),
            .I(N__5388));
    Span12Mux_h I__1260 (
            .O(N__5388),
            .I(N__5384));
    InMux I__1259 (
            .O(N__5387),
            .I(N__5381));
    Odrv12 I__1258 (
            .O(N__5384),
            .I(debouncedconsolereset));
    LocalMux I__1257 (
            .O(N__5381),
            .I(debouncedconsolereset));
    IoInMux I__1256 (
            .O(N__5376),
            .I(N__5373));
    LocalMux I__1255 (
            .O(N__5373),
            .I(\arse.apuresetoutregZ0 ));
    InMux I__1254 (
            .O(N__5370),
            .I(N__5365));
    InMux I__1253 (
            .O(N__5369),
            .I(N__5360));
    InMux I__1252 (
            .O(N__5368),
            .I(N__5360));
    LocalMux I__1251 (
            .O(N__5365),
            .I(arse_diveight_counter_1));
    LocalMux I__1250 (
            .O(N__5360),
            .I(arse_diveight_counter_1));
    InMux I__1249 (
            .O(N__5355),
            .I(N__5349));
    InMux I__1248 (
            .O(N__5354),
            .I(N__5346));
    InMux I__1247 (
            .O(N__5353),
            .I(N__5341));
    InMux I__1246 (
            .O(N__5352),
            .I(N__5341));
    LocalMux I__1245 (
            .O(N__5349),
            .I(arse_diveight_counter_0));
    LocalMux I__1244 (
            .O(N__5346),
            .I(arse_diveight_counter_0));
    LocalMux I__1243 (
            .O(N__5341),
            .I(arse_diveight_counter_0));
    CascadeMux I__1242 (
            .O(N__5334),
            .I(N__5331));
    InMux I__1241 (
            .O(N__5331),
            .I(N__5328));
    LocalMux I__1240 (
            .O(N__5328),
            .I(N__5322));
    InMux I__1239 (
            .O(N__5327),
            .I(N__5319));
    CascadeMux I__1238 (
            .O(N__5326),
            .I(N__5316));
    CascadeMux I__1237 (
            .O(N__5325),
            .I(N__5308));
    Span4Mux_v I__1236 (
            .O(N__5322),
            .I(N__5303));
    LocalMux I__1235 (
            .O(N__5319),
            .I(N__5303));
    InMux I__1234 (
            .O(N__5316),
            .I(N__5300));
    CascadeMux I__1233 (
            .O(N__5315),
            .I(N__5297));
    CascadeMux I__1232 (
            .O(N__5314),
            .I(N__5294));
    CascadeMux I__1231 (
            .O(N__5313),
            .I(N__5290));
    CascadeMux I__1230 (
            .O(N__5312),
            .I(N__5287));
    CascadeMux I__1229 (
            .O(N__5311),
            .I(N__5284));
    InMux I__1228 (
            .O(N__5308),
            .I(N__5279));
    Span4Mux_h I__1227 (
            .O(N__5303),
            .I(N__5274));
    LocalMux I__1226 (
            .O(N__5300),
            .I(N__5274));
    InMux I__1225 (
            .O(N__5297),
            .I(N__5271));
    InMux I__1224 (
            .O(N__5294),
            .I(N__5264));
    InMux I__1223 (
            .O(N__5293),
            .I(N__5264));
    InMux I__1222 (
            .O(N__5290),
            .I(N__5264));
    InMux I__1221 (
            .O(N__5287),
            .I(N__5259));
    InMux I__1220 (
            .O(N__5284),
            .I(N__5259));
    InMux I__1219 (
            .O(N__5283),
            .I(N__5256));
    InMux I__1218 (
            .O(N__5282),
            .I(N__5253));
    LocalMux I__1217 (
            .O(N__5279),
            .I(N__5250));
    Span4Mux_h I__1216 (
            .O(N__5274),
            .I(N__5247));
    LocalMux I__1215 (
            .O(N__5271),
            .I(N__5240));
    LocalMux I__1214 (
            .O(N__5264),
            .I(N__5240));
    LocalMux I__1213 (
            .O(N__5259),
            .I(N__5240));
    LocalMux I__1212 (
            .O(N__5256),
            .I(N__5235));
    LocalMux I__1211 (
            .O(N__5253),
            .I(N__5228));
    Span4Mux_v I__1210 (
            .O(N__5250),
            .I(N__5228));
    Span4Mux_v I__1209 (
            .O(N__5247),
            .I(N__5228));
    Span4Mux_v I__1208 (
            .O(N__5240),
            .I(N__5225));
    InMux I__1207 (
            .O(N__5239),
            .I(N__5220));
    InMux I__1206 (
            .O(N__5238),
            .I(N__5220));
    Span4Mux_h I__1205 (
            .O(N__5235),
            .I(N__5217));
    Odrv4 I__1204 (
            .O(N__5228),
            .I(delayConstantZ0Z_0));
    Odrv4 I__1203 (
            .O(N__5225),
            .I(delayConstantZ0Z_0));
    LocalMux I__1202 (
            .O(N__5220),
            .I(delayConstantZ0Z_0));
    Odrv4 I__1201 (
            .O(N__5217),
            .I(delayConstantZ0Z_0));
    InMux I__1200 (
            .O(N__5208),
            .I(N__5203));
    InMux I__1199 (
            .O(N__5207),
            .I(N__5200));
    InMux I__1198 (
            .O(N__5206),
            .I(N__5197));
    LocalMux I__1197 (
            .O(N__5203),
            .I(arse_diveight_counter_2));
    LocalMux I__1196 (
            .O(N__5200),
            .I(arse_diveight_counter_2));
    LocalMux I__1195 (
            .O(N__5197),
            .I(arse_diveight_counter_2));
    InMux I__1194 (
            .O(N__5190),
            .I(N__5187));
    LocalMux I__1193 (
            .O(N__5187),
            .I(\arse.diveight.doutZ0Z_1 ));
    SRMux I__1192 (
            .O(N__5184),
            .I(N__5181));
    LocalMux I__1191 (
            .O(N__5181),
            .I(N__5178));
    Odrv4 I__1190 (
            .O(N__5178),
            .I(\arse.diveight.cpuclkreset_i ));
    CascadeMux I__1189 (
            .O(N__5175),
            .I(\arse.m8_2_cascade_ ));
    InMux I__1188 (
            .O(N__5172),
            .I(N__5167));
    InMux I__1187 (
            .O(N__5171),
            .I(N__5162));
    InMux I__1186 (
            .O(N__5170),
            .I(N__5162));
    LocalMux I__1185 (
            .O(N__5167),
            .I(\arse.cpuresetcountZ0Z_0 ));
    LocalMux I__1184 (
            .O(N__5162),
            .I(\arse.cpuresetcountZ0Z_0 ));
    CascadeMux I__1183 (
            .O(N__5157),
            .I(N__5152));
    InMux I__1182 (
            .O(N__5156),
            .I(N__5149));
    InMux I__1181 (
            .O(N__5155),
            .I(N__5144));
    InMux I__1180 (
            .O(N__5152),
            .I(N__5144));
    LocalMux I__1179 (
            .O(N__5149),
            .I(\arse.cpuresetcountZ0Z_5 ));
    LocalMux I__1178 (
            .O(N__5144),
            .I(\arse.cpuresetcountZ0Z_5 ));
    CascadeMux I__1177 (
            .O(N__5139),
            .I(N__5135));
    InMux I__1176 (
            .O(N__5138),
            .I(N__5131));
    InMux I__1175 (
            .O(N__5135),
            .I(N__5126));
    InMux I__1174 (
            .O(N__5134),
            .I(N__5126));
    LocalMux I__1173 (
            .O(N__5131),
            .I(\arse.cpuresetcountZ0Z_1 ));
    LocalMux I__1172 (
            .O(N__5126),
            .I(\arse.cpuresetcountZ0Z_1 ));
    InMux I__1171 (
            .O(N__5121),
            .I(N__5116));
    InMux I__1170 (
            .O(N__5120),
            .I(N__5111));
    InMux I__1169 (
            .O(N__5119),
            .I(N__5111));
    LocalMux I__1168 (
            .O(N__5116),
            .I(\arse.cpuresetcountZ0Z_2 ));
    LocalMux I__1167 (
            .O(N__5111),
            .I(\arse.cpuresetcountZ0Z_2 ));
    CascadeMux I__1166 (
            .O(N__5106),
            .I(\arse.m12_2_cascade_ ));
    InMux I__1165 (
            .O(N__5103),
            .I(N__5098));
    InMux I__1164 (
            .O(N__5102),
            .I(N__5095));
    InMux I__1163 (
            .O(N__5101),
            .I(N__5092));
    LocalMux I__1162 (
            .O(N__5098),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1161 (
            .O(N__5095),
            .I(\arse.cpuresetcountZ0Z_4 ));
    LocalMux I__1160 (
            .O(N__5092),
            .I(\arse.cpuresetcountZ0Z_4 ));
    InMux I__1159 (
            .O(N__5085),
            .I(N__5082));
    LocalMux I__1158 (
            .O(N__5082),
            .I(\arse.cpuresetoutreg_1_sqmuxa ));
    InMux I__1157 (
            .O(N__5079),
            .I(N__5075));
    InMux I__1156 (
            .O(N__5078),
            .I(N__5072));
    LocalMux I__1155 (
            .O(N__5075),
            .I(\arse.cpuresetcountZ0Z_7 ));
    LocalMux I__1154 (
            .O(N__5072),
            .I(\arse.cpuresetcountZ0Z_7 ));
    InMux I__1153 (
            .O(N__5067),
            .I(N__5063));
    InMux I__1152 (
            .O(N__5066),
            .I(N__5060));
    LocalMux I__1151 (
            .O(N__5063),
            .I(\arse.cpuresetcountZ0Z_6 ));
    LocalMux I__1150 (
            .O(N__5060),
            .I(\arse.cpuresetcountZ0Z_6 ));
    InMux I__1149 (
            .O(N__5055),
            .I(N__5051));
    InMux I__1148 (
            .O(N__5054),
            .I(N__5048));
    LocalMux I__1147 (
            .O(N__5051),
            .I(\arse.cpuresetcountZ0Z_3 ));
    LocalMux I__1146 (
            .O(N__5048),
            .I(\arse.cpuresetcountZ0Z_3 ));
    InMux I__1145 (
            .O(N__5043),
            .I(N__5037));
    InMux I__1144 (
            .O(N__5042),
            .I(N__5037));
    LocalMux I__1143 (
            .O(N__5037),
            .I(\arse.m4_e_2 ));
    InMux I__1142 (
            .O(N__5034),
            .I(N__5031));
    LocalMux I__1141 (
            .O(N__5031),
            .I(\arse.cpuclkreset_1_sqmuxa ));
    SRMux I__1140 (
            .O(N__5028),
            .I(N__5023));
    SRMux I__1139 (
            .O(N__5027),
            .I(N__5020));
    SRMux I__1138 (
            .O(N__5026),
            .I(N__5017));
    LocalMux I__1137 (
            .O(N__5023),
            .I(N__5014));
    LocalMux I__1136 (
            .O(N__5020),
            .I(N__5011));
    LocalMux I__1135 (
            .O(N__5017),
            .I(N__5008));
    Span4Mux_v I__1134 (
            .O(N__5014),
            .I(N__5005));
    Odrv4 I__1133 (
            .O(N__5011),
            .I(debouncedconsolereset_i));
    Odrv4 I__1132 (
            .O(N__5008),
            .I(debouncedconsolereset_i));
    Odrv4 I__1131 (
            .O(N__5005),
            .I(debouncedconsolereset_i));
    InMux I__1130 (
            .O(N__4998),
            .I(N__4991));
    InMux I__1129 (
            .O(N__4997),
            .I(N__4987));
    InMux I__1128 (
            .O(N__4996),
            .I(N__4984));
    InMux I__1127 (
            .O(N__4995),
            .I(N__4981));
    CascadeMux I__1126 (
            .O(N__4994),
            .I(N__4978));
    LocalMux I__1125 (
            .O(N__4991),
            .I(N__4975));
    InMux I__1124 (
            .O(N__4990),
            .I(N__4972));
    LocalMux I__1123 (
            .O(N__4987),
            .I(N__4968));
    LocalMux I__1122 (
            .O(N__4984),
            .I(N__4965));
    LocalMux I__1121 (
            .O(N__4981),
            .I(N__4962));
    InMux I__1120 (
            .O(N__4978),
            .I(N__4959));
    Span4Mux_v I__1119 (
            .O(N__4975),
            .I(N__4956));
    LocalMux I__1118 (
            .O(N__4972),
            .I(N__4953));
    CascadeMux I__1117 (
            .O(N__4971),
            .I(N__4950));
    Sp12to4 I__1116 (
            .O(N__4968),
            .I(N__4941));
    Sp12to4 I__1115 (
            .O(N__4965),
            .I(N__4941));
    Sp12to4 I__1114 (
            .O(N__4962),
            .I(N__4941));
    LocalMux I__1113 (
            .O(N__4959),
            .I(N__4941));
    Span4Mux_h I__1112 (
            .O(N__4956),
            .I(N__4938));
    Span4Mux_v I__1111 (
            .O(N__4953),
            .I(N__4935));
    InMux I__1110 (
            .O(N__4950),
            .I(N__4932));
    Span12Mux_v I__1109 (
            .O(N__4941),
            .I(N__4929));
    Span4Mux_v I__1108 (
            .O(N__4938),
            .I(N__4926));
    Odrv4 I__1107 (
            .O(N__4935),
            .I(delayConstantZ0Z_3));
    LocalMux I__1106 (
            .O(N__4932),
            .I(delayConstantZ0Z_3));
    Odrv12 I__1105 (
            .O(N__4929),
            .I(delayConstantZ0Z_3));
    Odrv4 I__1104 (
            .O(N__4926),
            .I(delayConstantZ0Z_3));
    CascadeMux I__1103 (
            .O(N__4917),
            .I(arse_diveight_N_123_0_cascade_));
    InMux I__1102 (
            .O(N__4914),
            .I(\arse.un1_cpuresetcount_1_cry_1 ));
    InMux I__1101 (
            .O(N__4911),
            .I(\arse.un1_cpuresetcount_1_cry_2 ));
    InMux I__1100 (
            .O(N__4908),
            .I(\arse.un1_cpuresetcount_1_cry_3 ));
    InMux I__1099 (
            .O(N__4905),
            .I(\arse.un1_cpuresetcount_1_cry_4 ));
    InMux I__1098 (
            .O(N__4902),
            .I(\arse.un1_cpuresetcount_1_cry_5 ));
    InMux I__1097 (
            .O(N__4899),
            .I(\arse.un1_cpuresetcount_1_cry_6 ));
    IoInMux I__1096 (
            .O(N__4896),
            .I(N__4893));
    LocalMux I__1095 (
            .O(N__4893),
            .I(N__4889));
    InMux I__1094 (
            .O(N__4892),
            .I(N__4886));
    Span12Mux_s2_h I__1093 (
            .O(N__4889),
            .I(N__4883));
    LocalMux I__1092 (
            .O(N__4886),
            .I(\arse.cpuresetoutregZ0 ));
    Odrv12 I__1091 (
            .O(N__4883),
            .I(\arse.cpuresetoutregZ0 ));
    IoInMux I__1090 (
            .O(N__4878),
            .I(N__4875));
    LocalMux I__1089 (
            .O(N__4875),
            .I(N__4872));
    Span4Mux_s2_v I__1088 (
            .O(N__4872),
            .I(N__4868));
    InMux I__1087 (
            .O(N__4871),
            .I(N__4865));
    Span4Mux_h I__1086 (
            .O(N__4868),
            .I(N__4860));
    LocalMux I__1085 (
            .O(N__4865),
            .I(N__4857));
    CascadeMux I__1084 (
            .O(N__4864),
            .I(N__4854));
    InMux I__1083 (
            .O(N__4863),
            .I(N__4849));
    Span4Mux_h I__1082 (
            .O(N__4860),
            .I(N__4846));
    Sp12to4 I__1081 (
            .O(N__4857),
            .I(N__4843));
    InMux I__1080 (
            .O(N__4854),
            .I(N__4838));
    InMux I__1079 (
            .O(N__4853),
            .I(N__4838));
    InMux I__1078 (
            .O(N__4852),
            .I(N__4835));
    LocalMux I__1077 (
            .O(N__4849),
            .I(N__4831));
    Sp12to4 I__1076 (
            .O(N__4846),
            .I(N__4828));
    Span12Mux_v I__1075 (
            .O(N__4843),
            .I(N__4825));
    LocalMux I__1074 (
            .O(N__4838),
            .I(N__4822));
    LocalMux I__1073 (
            .O(N__4835),
            .I(N__4819));
    InMux I__1072 (
            .O(N__4834),
            .I(N__4816));
    Span4Mux_v I__1071 (
            .O(N__4831),
            .I(N__4813));
    Span12Mux_v I__1070 (
            .O(N__4828),
            .I(N__4810));
    Span12Mux_h I__1069 (
            .O(N__4825),
            .I(N__4807));
    Span12Mux_h I__1068 (
            .O(N__4822),
            .I(N__4802));
    Span12Mux_v I__1067 (
            .O(N__4819),
            .I(N__4802));
    LocalMux I__1066 (
            .O(N__4816),
            .I(N__4797));
    Sp12to4 I__1065 (
            .O(N__4813),
            .I(N__4797));
    Span12Mux_v I__1064 (
            .O(N__4810),
            .I(N__4792));
    Span12Mux_h I__1063 (
            .O(N__4807),
            .I(N__4792));
    Span12Mux_v I__1062 (
            .O(N__4802),
            .I(N__4789));
    Span12Mux_h I__1061 (
            .O(N__4797),
            .I(N__4786));
    Odrv12 I__1060 (
            .O(N__4792),
            .I(masterreset_c));
    Odrv12 I__1059 (
            .O(N__4789),
            .I(masterreset_c));
    Odrv12 I__1058 (
            .O(N__4786),
            .I(masterreset_c));
    CascadeMux I__1057 (
            .O(N__4779),
            .I(delayConstant17_i_cascade_));
    InMux I__1056 (
            .O(N__4776),
            .I(N__4773));
    LocalMux I__1055 (
            .O(N__4773),
            .I(un1_delayConstant_cry_0_c_RNOZ0));
    InMux I__1054 (
            .O(N__4770),
            .I(N__4767));
    LocalMux I__1053 (
            .O(N__4767),
            .I(olddn_RNIM5BH1Z0Z_4));
    InMux I__1052 (
            .O(N__4764),
            .I(N__4761));
    LocalMux I__1051 (
            .O(N__4761),
            .I(olddn_RNIM5BHZ0Z1));
    InMux I__1050 (
            .O(N__4758),
            .I(N__4755));
    LocalMux I__1049 (
            .O(N__4755),
            .I(N__4752));
    Span12Mux_v I__1048 (
            .O(N__4752),
            .I(N__4742));
    InMux I__1047 (
            .O(N__4751),
            .I(N__4739));
    InMux I__1046 (
            .O(N__4750),
            .I(N__4726));
    InMux I__1045 (
            .O(N__4749),
            .I(N__4726));
    InMux I__1044 (
            .O(N__4748),
            .I(N__4726));
    InMux I__1043 (
            .O(N__4747),
            .I(N__4726));
    InMux I__1042 (
            .O(N__4746),
            .I(N__4726));
    InMux I__1041 (
            .O(N__4745),
            .I(N__4726));
    Odrv12 I__1040 (
            .O(N__4742),
            .I(olddn_RNIEENHZ0));
    LocalMux I__1039 (
            .O(N__4739),
            .I(olddn_RNIEENHZ0));
    LocalMux I__1038 (
            .O(N__4726),
            .I(olddn_RNIEENHZ0));
    InMux I__1037 (
            .O(N__4719),
            .I(N__4716));
    LocalMux I__1036 (
            .O(N__4716),
            .I(N__4713));
    Span4Mux_h I__1035 (
            .O(N__4713),
            .I(N__4707));
    CascadeMux I__1034 (
            .O(N__4712),
            .I(N__4703));
    CascadeMux I__1033 (
            .O(N__4711),
            .I(N__4699));
    CascadeMux I__1032 (
            .O(N__4710),
            .I(N__4696));
    Span4Mux_v I__1031 (
            .O(N__4707),
            .I(N__4691));
    InMux I__1030 (
            .O(N__4706),
            .I(N__4688));
    InMux I__1029 (
            .O(N__4703),
            .I(N__4677));
    InMux I__1028 (
            .O(N__4702),
            .I(N__4677));
    InMux I__1027 (
            .O(N__4699),
            .I(N__4677));
    InMux I__1026 (
            .O(N__4696),
            .I(N__4677));
    InMux I__1025 (
            .O(N__4695),
            .I(N__4677));
    InMux I__1024 (
            .O(N__4694),
            .I(N__4674));
    Odrv4 I__1023 (
            .O(N__4691),
            .I(delayConstant17_i));
    LocalMux I__1022 (
            .O(N__4688),
            .I(delayConstant17_i));
    LocalMux I__1021 (
            .O(N__4677),
            .I(delayConstant17_i));
    LocalMux I__1020 (
            .O(N__4674),
            .I(delayConstant17_i));
    InMux I__1019 (
            .O(N__4665),
            .I(N__4662));
    LocalMux I__1018 (
            .O(N__4662),
            .I(olddn_RNIM5BH1Z0Z_2));
    InMux I__1017 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__1016 (
            .O(N__4656),
            .I(oldupZ0));
    InMux I__1015 (
            .O(N__4653),
            .I(N__4649));
    CascadeMux I__1014 (
            .O(N__4652),
            .I(N__4646));
    LocalMux I__1013 (
            .O(N__4649),
            .I(N__4643));
    InMux I__1012 (
            .O(N__4646),
            .I(N__4640));
    Span12Mux_s9_h I__1011 (
            .O(N__4643),
            .I(N__4637));
    LocalMux I__1010 (
            .O(N__4640),
            .I(\debounceup.counter19 ));
    Odrv12 I__1009 (
            .O(N__4637),
            .I(\debounceup.counter19 ));
    InMux I__1008 (
            .O(N__4632),
            .I(N__4629));
    LocalMux I__1007 (
            .O(N__4629),
            .I(N__4626));
    Span4Mux_v I__1006 (
            .O(N__4626),
            .I(N__4623));
    Sp12to4 I__1005 (
            .O(N__4623),
            .I(N__4620));
    Span12Mux_s6_h I__1004 (
            .O(N__4620),
            .I(N__4617));
    Odrv12 I__1003 (
            .O(N__4617),
            .I(delup_c));
    InMux I__1002 (
            .O(N__4614),
            .I(N__4610));
    InMux I__1001 (
            .O(N__4613),
            .I(N__4607));
    LocalMux I__1000 (
            .O(N__4610),
            .I(N__4588));
    LocalMux I__999 (
            .O(N__4607),
            .I(N__4585));
    CEMux I__998 (
            .O(N__4606),
            .I(N__4548));
    CEMux I__997 (
            .O(N__4605),
            .I(N__4548));
    CEMux I__996 (
            .O(N__4604),
            .I(N__4548));
    CEMux I__995 (
            .O(N__4603),
            .I(N__4548));
    CEMux I__994 (
            .O(N__4602),
            .I(N__4548));
    CEMux I__993 (
            .O(N__4601),
            .I(N__4548));
    CEMux I__992 (
            .O(N__4600),
            .I(N__4548));
    CEMux I__991 (
            .O(N__4599),
            .I(N__4548));
    CEMux I__990 (
            .O(N__4598),
            .I(N__4548));
    CEMux I__989 (
            .O(N__4597),
            .I(N__4548));
    CEMux I__988 (
            .O(N__4596),
            .I(N__4548));
    CEMux I__987 (
            .O(N__4595),
            .I(N__4548));
    CEMux I__986 (
            .O(N__4594),
            .I(N__4548));
    CEMux I__985 (
            .O(N__4593),
            .I(N__4548));
    CEMux I__984 (
            .O(N__4592),
            .I(N__4548));
    CEMux I__983 (
            .O(N__4591),
            .I(N__4548));
    Glb2LocalMux I__982 (
            .O(N__4588),
            .I(N__4548));
    Glb2LocalMux I__981 (
            .O(N__4585),
            .I(N__4548));
    GlobalMux I__980 (
            .O(N__4548),
            .I(N__4545));
    gio2CtrlBuf I__979 (
            .O(N__4545),
            .I(N_111_g));
    InMux I__978 (
            .O(N__4542),
            .I(N__4535));
    InMux I__977 (
            .O(N__4541),
            .I(N__4535));
    CascadeMux I__976 (
            .O(N__4540),
            .I(N__4532));
    LocalMux I__975 (
            .O(N__4535),
            .I(N__4529));
    InMux I__974 (
            .O(N__4532),
            .I(N__4526));
    Span12Mux_s10_v I__973 (
            .O(N__4529),
            .I(N__4523));
    LocalMux I__972 (
            .O(N__4526),
            .I(debouncedup));
    Odrv12 I__971 (
            .O(N__4523),
            .I(debouncedup));
    InMux I__970 (
            .O(N__4518),
            .I(N__4515));
    LocalMux I__969 (
            .O(N__4515),
            .I(N__4484));
    ClkMux I__968 (
            .O(N__4514),
            .I(N__4425));
    ClkMux I__967 (
            .O(N__4513),
            .I(N__4425));
    ClkMux I__966 (
            .O(N__4512),
            .I(N__4425));
    ClkMux I__965 (
            .O(N__4511),
            .I(N__4425));
    ClkMux I__964 (
            .O(N__4510),
            .I(N__4425));
    ClkMux I__963 (
            .O(N__4509),
            .I(N__4425));
    ClkMux I__962 (
            .O(N__4508),
            .I(N__4425));
    ClkMux I__961 (
            .O(N__4507),
            .I(N__4425));
    ClkMux I__960 (
            .O(N__4506),
            .I(N__4425));
    ClkMux I__959 (
            .O(N__4505),
            .I(N__4425));
    ClkMux I__958 (
            .O(N__4504),
            .I(N__4425));
    ClkMux I__957 (
            .O(N__4503),
            .I(N__4425));
    ClkMux I__956 (
            .O(N__4502),
            .I(N__4425));
    ClkMux I__955 (
            .O(N__4501),
            .I(N__4425));
    ClkMux I__954 (
            .O(N__4500),
            .I(N__4425));
    ClkMux I__953 (
            .O(N__4499),
            .I(N__4425));
    ClkMux I__952 (
            .O(N__4498),
            .I(N__4425));
    ClkMux I__951 (
            .O(N__4497),
            .I(N__4425));
    ClkMux I__950 (
            .O(N__4496),
            .I(N__4425));
    ClkMux I__949 (
            .O(N__4495),
            .I(N__4425));
    ClkMux I__948 (
            .O(N__4494),
            .I(N__4425));
    ClkMux I__947 (
            .O(N__4493),
            .I(N__4425));
    ClkMux I__946 (
            .O(N__4492),
            .I(N__4425));
    ClkMux I__945 (
            .O(N__4491),
            .I(N__4425));
    ClkMux I__944 (
            .O(N__4490),
            .I(N__4425));
    ClkMux I__943 (
            .O(N__4489),
            .I(N__4425));
    ClkMux I__942 (
            .O(N__4488),
            .I(N__4425));
    ClkMux I__941 (
            .O(N__4487),
            .I(N__4425));
    Glb2LocalMux I__940 (
            .O(N__4484),
            .I(N__4425));
    GlobalMux I__939 (
            .O(N__4425),
            .I(N__4422));
    gio2CtrlBuf I__938 (
            .O(N__4422),
            .I(PACKAGEPIN_0_c_g));
    InMux I__937 (
            .O(N__4419),
            .I(\arse.un1_cpuresetcount_1_cry_0 ));
    InMux I__936 (
            .O(N__4416),
            .I(N__4409));
    InMux I__935 (
            .O(N__4415),
            .I(N__4406));
    InMux I__934 (
            .O(N__4414),
            .I(N__4400));
    InMux I__933 (
            .O(N__4413),
            .I(N__4395));
    InMux I__932 (
            .O(N__4412),
            .I(N__4395));
    LocalMux I__931 (
            .O(N__4409),
            .I(N__4390));
    LocalMux I__930 (
            .O(N__4406),
            .I(N__4390));
    InMux I__929 (
            .O(N__4405),
            .I(N__4385));
    InMux I__928 (
            .O(N__4404),
            .I(N__4385));
    InMux I__927 (
            .O(N__4403),
            .I(N__4381));
    LocalMux I__926 (
            .O(N__4400),
            .I(N__4376));
    LocalMux I__925 (
            .O(N__4395),
            .I(N__4376));
    Span4Mux_v I__924 (
            .O(N__4390),
            .I(N__4369));
    LocalMux I__923 (
            .O(N__4385),
            .I(N__4369));
    InMux I__922 (
            .O(N__4384),
            .I(N__4366));
    LocalMux I__921 (
            .O(N__4381),
            .I(N__4363));
    Span4Mux_h I__920 (
            .O(N__4376),
            .I(N__4360));
    InMux I__919 (
            .O(N__4375),
            .I(N__4357));
    CascadeMux I__918 (
            .O(N__4374),
            .I(N__4354));
    Span4Mux_h I__917 (
            .O(N__4369),
            .I(N__4351));
    LocalMux I__916 (
            .O(N__4366),
            .I(N__4342));
    Sp12to4 I__915 (
            .O(N__4363),
            .I(N__4342));
    Sp12to4 I__914 (
            .O(N__4360),
            .I(N__4342));
    LocalMux I__913 (
            .O(N__4357),
            .I(N__4342));
    InMux I__912 (
            .O(N__4354),
            .I(N__4339));
    Span4Mux_v I__911 (
            .O(N__4351),
            .I(N__4336));
    Span12Mux_v I__910 (
            .O(N__4342),
            .I(N__4333));
    LocalMux I__909 (
            .O(N__4339),
            .I(delayConstantZ0Z_4));
    Odrv4 I__908 (
            .O(N__4336),
            .I(delayConstantZ0Z_4));
    Odrv12 I__907 (
            .O(N__4333),
            .I(delayConstantZ0Z_4));
    InMux I__906 (
            .O(N__4326),
            .I(un1_delayConstant_cry_3));
    InMux I__905 (
            .O(N__4323),
            .I(N__4318));
    CascadeMux I__904 (
            .O(N__4322),
            .I(N__4315));
    CascadeMux I__903 (
            .O(N__4321),
            .I(N__4312));
    LocalMux I__902 (
            .O(N__4318),
            .I(N__4308));
    InMux I__901 (
            .O(N__4315),
            .I(N__4305));
    InMux I__900 (
            .O(N__4312),
            .I(N__4300));
    CascadeMux I__899 (
            .O(N__4311),
            .I(N__4296));
    Span4Mux_v I__898 (
            .O(N__4308),
            .I(N__4289));
    LocalMux I__897 (
            .O(N__4305),
            .I(N__4289));
    CascadeMux I__896 (
            .O(N__4304),
            .I(N__4286));
    CascadeMux I__895 (
            .O(N__4303),
            .I(N__4282));
    LocalMux I__894 (
            .O(N__4300),
            .I(N__4279));
    InMux I__893 (
            .O(N__4299),
            .I(N__4274));
    InMux I__892 (
            .O(N__4296),
            .I(N__4274));
    CascadeMux I__891 (
            .O(N__4295),
            .I(N__4271));
    InMux I__890 (
            .O(N__4294),
            .I(N__4268));
    Span4Mux_v I__889 (
            .O(N__4289),
            .I(N__4265));
    InMux I__888 (
            .O(N__4286),
            .I(N__4260));
    InMux I__887 (
            .O(N__4285),
            .I(N__4260));
    InMux I__886 (
            .O(N__4282),
            .I(N__4256));
    Span4Mux_v I__885 (
            .O(N__4279),
            .I(N__4253));
    LocalMux I__884 (
            .O(N__4274),
            .I(N__4250));
    InMux I__883 (
            .O(N__4271),
            .I(N__4247));
    LocalMux I__882 (
            .O(N__4268),
            .I(N__4244));
    Span4Mux_h I__881 (
            .O(N__4265),
            .I(N__4239));
    LocalMux I__880 (
            .O(N__4260),
            .I(N__4239));
    CascadeMux I__879 (
            .O(N__4259),
            .I(N__4236));
    LocalMux I__878 (
            .O(N__4256),
            .I(N__4231));
    Sp12to4 I__877 (
            .O(N__4253),
            .I(N__4231));
    Sp12to4 I__876 (
            .O(N__4250),
            .I(N__4226));
    LocalMux I__875 (
            .O(N__4247),
            .I(N__4226));
    Span4Mux_v I__874 (
            .O(N__4244),
            .I(N__4223));
    Span4Mux_h I__873 (
            .O(N__4239),
            .I(N__4220));
    InMux I__872 (
            .O(N__4236),
            .I(N__4217));
    Span12Mux_h I__871 (
            .O(N__4231),
            .I(N__4214));
    Span12Mux_v I__870 (
            .O(N__4226),
            .I(N__4211));
    Span4Mux_h I__869 (
            .O(N__4223),
            .I(N__4206));
    Span4Mux_v I__868 (
            .O(N__4220),
            .I(N__4206));
    LocalMux I__867 (
            .O(N__4217),
            .I(delayConstantZ0Z_5));
    Odrv12 I__866 (
            .O(N__4214),
            .I(delayConstantZ0Z_5));
    Odrv12 I__865 (
            .O(N__4211),
            .I(delayConstantZ0Z_5));
    Odrv4 I__864 (
            .O(N__4206),
            .I(delayConstantZ0Z_5));
    InMux I__863 (
            .O(N__4197),
            .I(un1_delayConstant_cry_4));
    InMux I__862 (
            .O(N__4194),
            .I(N__4191));
    LocalMux I__861 (
            .O(N__4191),
            .I(N__4187));
    InMux I__860 (
            .O(N__4190),
            .I(N__4182));
    Span4Mux_h I__859 (
            .O(N__4187),
            .I(N__4178));
    InMux I__858 (
            .O(N__4186),
            .I(N__4175));
    InMux I__857 (
            .O(N__4185),
            .I(N__4172));
    LocalMux I__856 (
            .O(N__4182),
            .I(N__4168));
    InMux I__855 (
            .O(N__4181),
            .I(N__4165));
    Span4Mux_h I__854 (
            .O(N__4178),
            .I(N__4160));
    LocalMux I__853 (
            .O(N__4175),
            .I(N__4160));
    LocalMux I__852 (
            .O(N__4172),
            .I(N__4157));
    CascadeMux I__851 (
            .O(N__4171),
            .I(N__4154));
    Sp12to4 I__850 (
            .O(N__4168),
            .I(N__4149));
    LocalMux I__849 (
            .O(N__4165),
            .I(N__4149));
    Span4Mux_h I__848 (
            .O(N__4160),
            .I(N__4146));
    Span12Mux_h I__847 (
            .O(N__4157),
            .I(N__4143));
    InMux I__846 (
            .O(N__4154),
            .I(N__4140));
    Span12Mux_v I__845 (
            .O(N__4149),
            .I(N__4137));
    Span4Mux_v I__844 (
            .O(N__4146),
            .I(N__4134));
    Odrv12 I__843 (
            .O(N__4143),
            .I(delayConstantZ0Z_6));
    LocalMux I__842 (
            .O(N__4140),
            .I(delayConstantZ0Z_6));
    Odrv12 I__841 (
            .O(N__4137),
            .I(delayConstantZ0Z_6));
    Odrv4 I__840 (
            .O(N__4134),
            .I(delayConstantZ0Z_6));
    InMux I__839 (
            .O(N__4125),
            .I(un1_delayConstant_cry_5));
    InMux I__838 (
            .O(N__4122),
            .I(un1_delayConstant_cry_6));
    InMux I__837 (
            .O(N__4119),
            .I(N__4115));
    CascadeMux I__836 (
            .O(N__4118),
            .I(N__4111));
    LocalMux I__835 (
            .O(N__4115),
            .I(N__4106));
    InMux I__834 (
            .O(N__4114),
            .I(N__4101));
    InMux I__833 (
            .O(N__4111),
            .I(N__4101));
    CascadeMux I__832 (
            .O(N__4110),
            .I(N__4098));
    InMux I__831 (
            .O(N__4109),
            .I(N__4095));
    Span4Mux_h I__830 (
            .O(N__4106),
            .I(N__4090));
    LocalMux I__829 (
            .O(N__4101),
            .I(N__4090));
    InMux I__828 (
            .O(N__4098),
            .I(N__4086));
    LocalMux I__827 (
            .O(N__4095),
            .I(N__4083));
    Span4Mux_v I__826 (
            .O(N__4090),
            .I(N__4080));
    CascadeMux I__825 (
            .O(N__4089),
            .I(N__4077));
    LocalMux I__824 (
            .O(N__4086),
            .I(N__4074));
    Span4Mux_v I__823 (
            .O(N__4083),
            .I(N__4069));
    Span4Mux_h I__822 (
            .O(N__4080),
            .I(N__4069));
    InMux I__821 (
            .O(N__4077),
            .I(N__4066));
    Span12Mux_h I__820 (
            .O(N__4074),
            .I(N__4063));
    Span4Mux_v I__819 (
            .O(N__4069),
            .I(N__4060));
    LocalMux I__818 (
            .O(N__4066),
            .I(delayConstantZ0Z_7));
    Odrv12 I__817 (
            .O(N__4063),
            .I(delayConstantZ0Z_7));
    Odrv4 I__816 (
            .O(N__4060),
            .I(delayConstantZ0Z_7));
    SRMux I__815 (
            .O(N__4053),
            .I(N__4035));
    SRMux I__814 (
            .O(N__4052),
            .I(N__4035));
    SRMux I__813 (
            .O(N__4051),
            .I(N__4035));
    SRMux I__812 (
            .O(N__4050),
            .I(N__4035));
    SRMux I__811 (
            .O(N__4049),
            .I(N__4035));
    SRMux I__810 (
            .O(N__4048),
            .I(N__4035));
    GlobalMux I__809 (
            .O(N__4035),
            .I(N__4032));
    gio2CtrlBuf I__808 (
            .O(N__4032),
            .I(masterreset_c_i_g));
    InMux I__807 (
            .O(N__4029),
            .I(N__4026));
    LocalMux I__806 (
            .O(N__4026),
            .I(olddnZ0));
    CascadeMux I__805 (
            .O(N__4023),
            .I(N__4020));
    InMux I__804 (
            .O(N__4020),
            .I(N__4015));
    InMux I__803 (
            .O(N__4019),
            .I(N__4010));
    InMux I__802 (
            .O(N__4018),
            .I(N__4010));
    LocalMux I__801 (
            .O(N__4015),
            .I(debounceddn));
    LocalMux I__800 (
            .O(N__4010),
            .I(debounceddn));
    CascadeMux I__799 (
            .O(N__4005),
            .I(olddn_RNIEENHZ0_cascade_));
    InMux I__798 (
            .O(N__4002),
            .I(N__3999));
    LocalMux I__797 (
            .O(N__3999),
            .I(olddn_RNIM5BH1Z0Z_0));
    InMux I__796 (
            .O(N__3996),
            .I(N__3993));
    LocalMux I__795 (
            .O(N__3993),
            .I(olddn_RNIM5BH1Z0Z_3));
    InMux I__794 (
            .O(N__3990),
            .I(N__3987));
    LocalMux I__793 (
            .O(N__3987),
            .I(olddn_RNIM5BH1Z0Z_1));
    CascadeMux I__792 (
            .O(N__3984),
            .I(N__3981));
    InMux I__791 (
            .O(N__3981),
            .I(N__3976));
    InMux I__790 (
            .O(N__3980),
            .I(N__3973));
    InMux I__789 (
            .O(N__3979),
            .I(N__3970));
    LocalMux I__788 (
            .O(N__3976),
            .I(N__3965));
    LocalMux I__787 (
            .O(N__3973),
            .I(N__3965));
    LocalMux I__786 (
            .O(N__3970),
            .I(\debouncedn.counter19_2 ));
    Odrv4 I__785 (
            .O(N__3965),
            .I(\debouncedn.counter19_2 ));
    InMux I__784 (
            .O(N__3960),
            .I(\debouncedn.un3_counter_1_cry_3 ));
    InMux I__783 (
            .O(N__3957),
            .I(N__3951));
    InMux I__782 (
            .O(N__3956),
            .I(N__3948));
    InMux I__781 (
            .O(N__3955),
            .I(N__3945));
    InMux I__780 (
            .O(N__3954),
            .I(N__3942));
    LocalMux I__779 (
            .O(N__3951),
            .I(\debouncedn.counterZ0Z_4 ));
    LocalMux I__778 (
            .O(N__3948),
            .I(\debouncedn.counterZ0Z_4 ));
    LocalMux I__777 (
            .O(N__3945),
            .I(\debouncedn.counterZ0Z_4 ));
    LocalMux I__776 (
            .O(N__3942),
            .I(\debouncedn.counterZ0Z_4 ));
    InMux I__775 (
            .O(N__3933),
            .I(N__3927));
    CascadeMux I__774 (
            .O(N__3932),
            .I(N__3924));
    InMux I__773 (
            .O(N__3931),
            .I(N__3921));
    InMux I__772 (
            .O(N__3930),
            .I(N__3918));
    LocalMux I__771 (
            .O(N__3927),
            .I(N__3915));
    InMux I__770 (
            .O(N__3924),
            .I(N__3912));
    LocalMux I__769 (
            .O(N__3921),
            .I(\debouncedn.counterZ0Z_0 ));
    LocalMux I__768 (
            .O(N__3918),
            .I(\debouncedn.counterZ0Z_0 ));
    Odrv4 I__767 (
            .O(N__3915),
            .I(\debouncedn.counterZ0Z_0 ));
    LocalMux I__766 (
            .O(N__3912),
            .I(\debouncedn.counterZ0Z_0 ));
    InMux I__765 (
            .O(N__3903),
            .I(N__3899));
    InMux I__764 (
            .O(N__3902),
            .I(N__3895));
    LocalMux I__763 (
            .O(N__3899),
            .I(N__3892));
    InMux I__762 (
            .O(N__3898),
            .I(N__3889));
    LocalMux I__761 (
            .O(N__3895),
            .I(\debouncedn.counterZ0Z_1 ));
    Odrv4 I__760 (
            .O(N__3892),
            .I(\debouncedn.counterZ0Z_1 ));
    LocalMux I__759 (
            .O(N__3889),
            .I(\debouncedn.counterZ0Z_1 ));
    InMux I__758 (
            .O(N__3882),
            .I(N__3879));
    LocalMux I__757 (
            .O(N__3879),
            .I(N__3875));
    InMux I__756 (
            .O(N__3878),
            .I(N__3872));
    Span4Mux_h I__755 (
            .O(N__3875),
            .I(N__3869));
    LocalMux I__754 (
            .O(N__3872),
            .I(\debouncedn.counter19 ));
    Odrv4 I__753 (
            .O(N__3869),
            .I(\debouncedn.counter19 ));
    InMux I__752 (
            .O(N__3864),
            .I(N__3861));
    LocalMux I__751 (
            .O(N__3861),
            .I(N__3858));
    Span4Mux_v I__750 (
            .O(N__3858),
            .I(N__3855));
    Span4Mux_h I__749 (
            .O(N__3855),
            .I(N__3852));
    Sp12to4 I__748 (
            .O(N__3852),
            .I(N__3849));
    Span12Mux_h I__747 (
            .O(N__3849),
            .I(N__3846));
    Span12Mux_v I__746 (
            .O(N__3846),
            .I(N__3843));
    Odrv12 I__745 (
            .O(N__3843),
            .I(deldn_c));
    IoInMux I__744 (
            .O(N__3840),
            .I(N__3837));
    LocalMux I__743 (
            .O(N__3837),
            .I(N__3833));
    IoInMux I__742 (
            .O(N__3836),
            .I(N__3829));
    IoSpan4Mux I__741 (
            .O(N__3833),
            .I(N__3826));
    IoInMux I__740 (
            .O(N__3832),
            .I(N__3823));
    LocalMux I__739 (
            .O(N__3829),
            .I(N__3820));
    IoSpan4Mux I__738 (
            .O(N__3826),
            .I(N__3814));
    LocalMux I__737 (
            .O(N__3823),
            .I(N__3814));
    IoSpan4Mux I__736 (
            .O(N__3820),
            .I(N__3811));
    IoInMux I__735 (
            .O(N__3819),
            .I(N__3808));
    IoSpan4Mux I__734 (
            .O(N__3814),
            .I(N__3805));
    IoSpan4Mux I__733 (
            .O(N__3811),
            .I(N__3800));
    LocalMux I__732 (
            .O(N__3808),
            .I(N__3800));
    Span4Mux_s0_h I__731 (
            .O(N__3805),
            .I(N__3797));
    IoSpan4Mux I__730 (
            .O(N__3800),
            .I(N__3794));
    Sp12to4 I__729 (
            .O(N__3797),
            .I(N__3791));
    Span4Mux_s3_v I__728 (
            .O(N__3794),
            .I(N__3788));
    Span12Mux_v I__727 (
            .O(N__3791),
            .I(N__3785));
    Span4Mux_v I__726 (
            .O(N__3788),
            .I(N__3782));
    Odrv12 I__725 (
            .O(N__3785),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__724 (
            .O(N__3782),
            .I(CONSTANT_ONE_NET));
    InMux I__723 (
            .O(N__3777),
            .I(un1_delayConstant_cry_0));
    InMux I__722 (
            .O(N__3774),
            .I(un1_delayConstant_cry_1));
    InMux I__721 (
            .O(N__3771),
            .I(un1_delayConstant_cry_2));
    IoInMux I__720 (
            .O(N__3768),
            .I(N__3765));
    LocalMux I__719 (
            .O(N__3765),
            .I(N__3762));
    Span4Mux_s2_v I__718 (
            .O(N__3762),
            .I(N__3759));
    Span4Mux_h I__717 (
            .O(N__3759),
            .I(N__3756));
    Odrv4 I__716 (
            .O(N__3756),
            .I(lcol1_c));
    InMux I__715 (
            .O(N__3753),
            .I(N__3749));
    InMux I__714 (
            .O(N__3752),
            .I(N__3746));
    LocalMux I__713 (
            .O(N__3749),
            .I(N__3740));
    LocalMux I__712 (
            .O(N__3746),
            .I(N__3740));
    CascadeMux I__711 (
            .O(N__3745),
            .I(N__3733));
    Span4Mux_v I__710 (
            .O(N__3740),
            .I(N__3729));
    InMux I__709 (
            .O(N__3739),
            .I(N__3726));
    CascadeMux I__708 (
            .O(N__3738),
            .I(N__3722));
    InMux I__707 (
            .O(N__3737),
            .I(N__3716));
    InMux I__706 (
            .O(N__3736),
            .I(N__3711));
    InMux I__705 (
            .O(N__3733),
            .I(N__3711));
    InMux I__704 (
            .O(N__3732),
            .I(N__3706));
    Sp12to4 I__703 (
            .O(N__3729),
            .I(N__3701));
    LocalMux I__702 (
            .O(N__3726),
            .I(N__3701));
    InMux I__701 (
            .O(N__3725),
            .I(N__3698));
    InMux I__700 (
            .O(N__3722),
            .I(N__3693));
    InMux I__699 (
            .O(N__3721),
            .I(N__3693));
    CascadeMux I__698 (
            .O(N__3720),
            .I(N__3688));
    InMux I__697 (
            .O(N__3719),
            .I(N__3683));
    LocalMux I__696 (
            .O(N__3716),
            .I(N__3678));
    LocalMux I__695 (
            .O(N__3711),
            .I(N__3678));
    InMux I__694 (
            .O(N__3710),
            .I(N__3673));
    InMux I__693 (
            .O(N__3709),
            .I(N__3673));
    LocalMux I__692 (
            .O(N__3706),
            .I(N__3667));
    Span12Mux_h I__691 (
            .O(N__3701),
            .I(N__3667));
    LocalMux I__690 (
            .O(N__3698),
            .I(N__3661));
    LocalMux I__689 (
            .O(N__3693),
            .I(N__3661));
    InMux I__688 (
            .O(N__3692),
            .I(N__3654));
    InMux I__687 (
            .O(N__3691),
            .I(N__3645));
    InMux I__686 (
            .O(N__3688),
            .I(N__3645));
    InMux I__685 (
            .O(N__3687),
            .I(N__3645));
    InMux I__684 (
            .O(N__3686),
            .I(N__3645));
    LocalMux I__683 (
            .O(N__3683),
            .I(N__3638));
    Span4Mux_v I__682 (
            .O(N__3678),
            .I(N__3638));
    LocalMux I__681 (
            .O(N__3673),
            .I(N__3638));
    InMux I__680 (
            .O(N__3672),
            .I(N__3635));
    Span12Mux_v I__679 (
            .O(N__3667),
            .I(N__3632));
    InMux I__678 (
            .O(N__3666),
            .I(N__3629));
    Span4Mux_v I__677 (
            .O(N__3661),
            .I(N__3626));
    InMux I__676 (
            .O(N__3660),
            .I(N__3621));
    InMux I__675 (
            .O(N__3659),
            .I(N__3621));
    InMux I__674 (
            .O(N__3658),
            .I(N__3616));
    InMux I__673 (
            .O(N__3657),
            .I(N__3616));
    LocalMux I__672 (
            .O(N__3654),
            .I(N__3613));
    LocalMux I__671 (
            .O(N__3645),
            .I(N__3608));
    Span4Mux_h I__670 (
            .O(N__3638),
            .I(N__3608));
    LocalMux I__669 (
            .O(N__3635),
            .I(colZ0Z_1));
    Odrv12 I__668 (
            .O(N__3632),
            .I(colZ0Z_1));
    LocalMux I__667 (
            .O(N__3629),
            .I(colZ0Z_1));
    Odrv4 I__666 (
            .O(N__3626),
            .I(colZ0Z_1));
    LocalMux I__665 (
            .O(N__3621),
            .I(colZ0Z_1));
    LocalMux I__664 (
            .O(N__3616),
            .I(colZ0Z_1));
    Odrv4 I__663 (
            .O(N__3613),
            .I(colZ0Z_1));
    Odrv4 I__662 (
            .O(N__3608),
            .I(colZ0Z_1));
    InMux I__661 (
            .O(N__3591),
            .I(N__3588));
    LocalMux I__660 (
            .O(N__3588),
            .I(N__3583));
    CascadeMux I__659 (
            .O(N__3587),
            .I(N__3576));
    CascadeMux I__658 (
            .O(N__3586),
            .I(N__3573));
    Span4Mux_h I__657 (
            .O(N__3583),
            .I(N__3568));
    InMux I__656 (
            .O(N__3582),
            .I(N__3565));
    InMux I__655 (
            .O(N__3581),
            .I(N__3562));
    CascadeMux I__654 (
            .O(N__3580),
            .I(N__3549));
    InMux I__653 (
            .O(N__3579),
            .I(N__3546));
    InMux I__652 (
            .O(N__3576),
            .I(N__3541));
    InMux I__651 (
            .O(N__3573),
            .I(N__3541));
    InMux I__650 (
            .O(N__3572),
            .I(N__3538));
    InMux I__649 (
            .O(N__3571),
            .I(N__3535));
    Span4Mux_h I__648 (
            .O(N__3568),
            .I(N__3532));
    LocalMux I__647 (
            .O(N__3565),
            .I(N__3529));
    LocalMux I__646 (
            .O(N__3562),
            .I(N__3526));
    InMux I__645 (
            .O(N__3561),
            .I(N__3517));
    InMux I__644 (
            .O(N__3560),
            .I(N__3517));
    InMux I__643 (
            .O(N__3559),
            .I(N__3517));
    InMux I__642 (
            .O(N__3558),
            .I(N__3517));
    InMux I__641 (
            .O(N__3557),
            .I(N__3514));
    InMux I__640 (
            .O(N__3556),
            .I(N__3509));
    InMux I__639 (
            .O(N__3555),
            .I(N__3509));
    InMux I__638 (
            .O(N__3554),
            .I(N__3505));
    InMux I__637 (
            .O(N__3553),
            .I(N__3500));
    InMux I__636 (
            .O(N__3552),
            .I(N__3500));
    InMux I__635 (
            .O(N__3549),
            .I(N__3497));
    LocalMux I__634 (
            .O(N__3546),
            .I(N__3492));
    LocalMux I__633 (
            .O(N__3541),
            .I(N__3492));
    LocalMux I__632 (
            .O(N__3538),
            .I(N__3489));
    LocalMux I__631 (
            .O(N__3535),
            .I(N__3479));
    Sp12to4 I__630 (
            .O(N__3532),
            .I(N__3479));
    Span12Mux_h I__629 (
            .O(N__3529),
            .I(N__3479));
    Sp12to4 I__628 (
            .O(N__3526),
            .I(N__3479));
    LocalMux I__627 (
            .O(N__3517),
            .I(N__3469));
    LocalMux I__626 (
            .O(N__3514),
            .I(N__3469));
    LocalMux I__625 (
            .O(N__3509),
            .I(N__3466));
    InMux I__624 (
            .O(N__3508),
            .I(N__3463));
    LocalMux I__623 (
            .O(N__3505),
            .I(N__3458));
    LocalMux I__622 (
            .O(N__3500),
            .I(N__3458));
    LocalMux I__621 (
            .O(N__3497),
            .I(N__3453));
    Span4Mux_h I__620 (
            .O(N__3492),
            .I(N__3453));
    Span4Mux_h I__619 (
            .O(N__3489),
            .I(N__3450));
    InMux I__618 (
            .O(N__3488),
            .I(N__3447));
    Span12Mux_v I__617 (
            .O(N__3479),
            .I(N__3444));
    InMux I__616 (
            .O(N__3478),
            .I(N__3437));
    InMux I__615 (
            .O(N__3477),
            .I(N__3437));
    InMux I__614 (
            .O(N__3476),
            .I(N__3437));
    InMux I__613 (
            .O(N__3475),
            .I(N__3432));
    InMux I__612 (
            .O(N__3474),
            .I(N__3432));
    Span4Mux_v I__611 (
            .O(N__3469),
            .I(N__3427));
    Span4Mux_h I__610 (
            .O(N__3466),
            .I(N__3427));
    LocalMux I__609 (
            .O(N__3463),
            .I(N__3420));
    Span4Mux_v I__608 (
            .O(N__3458),
            .I(N__3420));
    Span4Mux_v I__607 (
            .O(N__3453),
            .I(N__3420));
    Odrv4 I__606 (
            .O(N__3450),
            .I(colZ0Z_0));
    LocalMux I__605 (
            .O(N__3447),
            .I(colZ0Z_0));
    Odrv12 I__604 (
            .O(N__3444),
            .I(colZ0Z_0));
    LocalMux I__603 (
            .O(N__3437),
            .I(colZ0Z_0));
    LocalMux I__602 (
            .O(N__3432),
            .I(colZ0Z_0));
    Odrv4 I__601 (
            .O(N__3427),
            .I(colZ0Z_0));
    Odrv4 I__600 (
            .O(N__3420),
            .I(colZ0Z_0));
    IoInMux I__599 (
            .O(N__3405),
            .I(N__3402));
    LocalMux I__598 (
            .O(N__3402),
            .I(N__3399));
    IoSpan4Mux I__597 (
            .O(N__3399),
            .I(N__3396));
    Odrv4 I__596 (
            .O(N__3396),
            .I(lcol2_c));
    CascadeMux I__595 (
            .O(N__3393),
            .I(\debouncedn.counter19_2_cascade_ ));
    CascadeMux I__594 (
            .O(N__3390),
            .I(\debouncedn.counter19_cascade_ ));
    InMux I__593 (
            .O(N__3387),
            .I(N__3383));
    InMux I__592 (
            .O(N__3386),
            .I(N__3380));
    LocalMux I__591 (
            .O(N__3383),
            .I(\debouncedn.counterZ0Z_2 ));
    LocalMux I__590 (
            .O(N__3380),
            .I(\debouncedn.counterZ0Z_2 ));
    InMux I__589 (
            .O(N__3375),
            .I(N__3372));
    LocalMux I__588 (
            .O(N__3372),
            .I(\debouncedn.counter_RNO_0_1_2 ));
    InMux I__587 (
            .O(N__3369),
            .I(\debouncedn.un3_counter_1_cry_1 ));
    InMux I__586 (
            .O(N__3366),
            .I(N__3362));
    InMux I__585 (
            .O(N__3365),
            .I(N__3359));
    LocalMux I__584 (
            .O(N__3362),
            .I(\debouncedn.counterZ0Z_3 ));
    LocalMux I__583 (
            .O(N__3359),
            .I(\debouncedn.counterZ0Z_3 ));
    InMux I__582 (
            .O(N__3354),
            .I(\debouncedn.un3_counter_1_cry_2 ));
    InMux I__581 (
            .O(N__3351),
            .I(N__3348));
    LocalMux I__580 (
            .O(N__3348),
            .I(N__3344));
    CascadeMux I__579 (
            .O(N__3347),
            .I(N__3339));
    Span12Mux_v I__578 (
            .O(N__3344),
            .I(N__3336));
    InMux I__577 (
            .O(N__3343),
            .I(N__3331));
    InMux I__576 (
            .O(N__3342),
            .I(N__3331));
    InMux I__575 (
            .O(N__3339),
            .I(N__3328));
    Odrv12 I__574 (
            .O(N__3336),
            .I(\debounceup.counterZ0Z_0 ));
    LocalMux I__573 (
            .O(N__3331),
            .I(\debounceup.counterZ0Z_0 ));
    LocalMux I__572 (
            .O(N__3328),
            .I(\debounceup.counterZ0Z_0 ));
    InMux I__571 (
            .O(N__3321),
            .I(N__3317));
    InMux I__570 (
            .O(N__3320),
            .I(N__3314));
    LocalMux I__569 (
            .O(N__3317),
            .I(N__3308));
    LocalMux I__568 (
            .O(N__3314),
            .I(N__3308));
    InMux I__567 (
            .O(N__3313),
            .I(N__3305));
    Span4Mux_v I__566 (
            .O(N__3308),
            .I(N__3302));
    LocalMux I__565 (
            .O(N__3305),
            .I(N__3297));
    Span4Mux_h I__564 (
            .O(N__3302),
            .I(N__3297));
    Odrv4 I__563 (
            .O(N__3297),
            .I(\debounceup.counterZ0Z_1 ));
    InMux I__562 (
            .O(N__3294),
            .I(N__3291));
    LocalMux I__561 (
            .O(N__3291),
            .I(\dig2.m49_bm ));
    InMux I__560 (
            .O(N__3288),
            .I(N__3285));
    LocalMux I__559 (
            .O(N__3285),
            .I(\dig2.m49_am ));
    InMux I__558 (
            .O(N__3282),
            .I(N__3279));
    LocalMux I__557 (
            .O(N__3279),
            .I(\dig2.m33_am ));
    CascadeMux I__556 (
            .O(N__3276),
            .I(\dig2.m33_bm_cascade_ ));
    IoInMux I__555 (
            .O(N__3273),
            .I(N__3270));
    LocalMux I__554 (
            .O(N__3270),
            .I(N__3267));
    Span12Mux_s4_v I__553 (
            .O(N__3267),
            .I(N__3264));
    Span12Mux_v I__552 (
            .O(N__3264),
            .I(N__3261));
    Span12Mux_h I__551 (
            .O(N__3261),
            .I(N__3258));
    Odrv12 I__550 (
            .O(N__3258),
            .I(leds_1_i_2));
    CascadeMux I__549 (
            .O(N__3255),
            .I(\dig2.N_25_cascade_ ));
    InMux I__548 (
            .O(N__3252),
            .I(N__3249));
    LocalMux I__547 (
            .O(N__3249),
            .I(\dig2.leds_17_i_0_ns_1_2 ));
    InMux I__546 (
            .O(N__3246),
            .I(N__3243));
    LocalMux I__545 (
            .O(N__3243),
            .I(\dig2.i2_mux ));
    InMux I__544 (
            .O(N__3240),
            .I(N__3237));
    LocalMux I__543 (
            .O(N__3237),
            .I(\debounceconsolereset.counter_RNO_0Z0Z_2 ));
    InMux I__542 (
            .O(N__3234),
            .I(\debounceconsolereset.un3_counter_1_cry_1 ));
    InMux I__541 (
            .O(N__3231),
            .I(\debounceconsolereset.un3_counter_1_cry_2 ));
    InMux I__540 (
            .O(N__3228),
            .I(\debounceconsolereset.un3_counter_1_cry_3 ));
    InMux I__539 (
            .O(N__3225),
            .I(N__3221));
    InMux I__538 (
            .O(N__3224),
            .I(N__3218));
    LocalMux I__537 (
            .O(N__3221),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    LocalMux I__536 (
            .O(N__3218),
            .I(\debounceconsolereset.counterZ0Z_3 ));
    InMux I__535 (
            .O(N__3213),
            .I(N__3209));
    InMux I__534 (
            .O(N__3212),
            .I(N__3206));
    LocalMux I__533 (
            .O(N__3209),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    LocalMux I__532 (
            .O(N__3206),
            .I(\debounceconsolereset.counterZ0Z_2 ));
    CascadeMux I__531 (
            .O(N__3201),
            .I(N__3197));
    InMux I__530 (
            .O(N__3200),
            .I(N__3193));
    InMux I__529 (
            .O(N__3197),
            .I(N__3188));
    InMux I__528 (
            .O(N__3196),
            .I(N__3188));
    LocalMux I__527 (
            .O(N__3193),
            .I(\debounceconsolereset.counter19_2 ));
    LocalMux I__526 (
            .O(N__3188),
            .I(\debounceconsolereset.counter19_2 ));
    InMux I__525 (
            .O(N__3183),
            .I(N__3175));
    InMux I__524 (
            .O(N__3182),
            .I(N__3175));
    InMux I__523 (
            .O(N__3181),
            .I(N__3172));
    InMux I__522 (
            .O(N__3180),
            .I(N__3169));
    LocalMux I__521 (
            .O(N__3175),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    LocalMux I__520 (
            .O(N__3172),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    LocalMux I__519 (
            .O(N__3169),
            .I(\debounceconsolereset.counterZ0Z_4 ));
    CascadeMux I__518 (
            .O(N__3162),
            .I(N__3158));
    InMux I__517 (
            .O(N__3161),
            .I(N__3154));
    InMux I__516 (
            .O(N__3158),
            .I(N__3151));
    InMux I__515 (
            .O(N__3157),
            .I(N__3148));
    LocalMux I__514 (
            .O(N__3154),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    LocalMux I__513 (
            .O(N__3151),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    LocalMux I__512 (
            .O(N__3148),
            .I(\debounceconsolereset.counterZ0Z_1 ));
    CascadeMux I__511 (
            .O(N__3141),
            .I(\debounceconsolereset.counter19_2_cascade_ ));
    InMux I__510 (
            .O(N__3138),
            .I(N__3130));
    InMux I__509 (
            .O(N__3137),
            .I(N__3130));
    InMux I__508 (
            .O(N__3136),
            .I(N__3127));
    InMux I__507 (
            .O(N__3135),
            .I(N__3124));
    LocalMux I__506 (
            .O(N__3130),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    LocalMux I__505 (
            .O(N__3127),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    LocalMux I__504 (
            .O(N__3124),
            .I(\debounceconsolereset.counterZ0Z_0 ));
    CascadeMux I__503 (
            .O(N__3117),
            .I(N__3114));
    InMux I__502 (
            .O(N__3114),
            .I(N__3109));
    InMux I__501 (
            .O(N__3113),
            .I(N__3106));
    InMux I__500 (
            .O(N__3112),
            .I(N__3103));
    LocalMux I__499 (
            .O(N__3109),
            .I(\debounceconsolereset.counter19 ));
    LocalMux I__498 (
            .O(N__3106),
            .I(\debounceconsolereset.counter19 ));
    LocalMux I__497 (
            .O(N__3103),
            .I(\debounceconsolereset.counter19 ));
    CascadeMux I__496 (
            .O(N__3096),
            .I(N__3092));
    InMux I__495 (
            .O(N__3095),
            .I(N__3088));
    InMux I__494 (
            .O(N__3092),
            .I(N__3083));
    InMux I__493 (
            .O(N__3091),
            .I(N__3080));
    LocalMux I__492 (
            .O(N__3088),
            .I(N__3077));
    InMux I__491 (
            .O(N__3087),
            .I(N__3074));
    InMux I__490 (
            .O(N__3086),
            .I(N__3071));
    LocalMux I__489 (
            .O(N__3083),
            .I(N__3068));
    LocalMux I__488 (
            .O(N__3080),
            .I(col_1_1));
    Odrv4 I__487 (
            .O(N__3077),
            .I(col_1_1));
    LocalMux I__486 (
            .O(N__3074),
            .I(col_1_1));
    LocalMux I__485 (
            .O(N__3071),
            .I(col_1_1));
    Odrv12 I__484 (
            .O(N__3068),
            .I(col_1_1));
    InMux I__483 (
            .O(N__3057),
            .I(N__3054));
    LocalMux I__482 (
            .O(N__3054),
            .I(N__3051));
    Odrv4 I__481 (
            .O(N__3051),
            .I(\dig2.m54_bm ));
    InMux I__480 (
            .O(N__3048),
            .I(N__3045));
    LocalMux I__479 (
            .O(N__3045),
            .I(N__3042));
    Odrv4 I__478 (
            .O(N__3042),
            .I(\dig2.leds_17_i_ns_1_1 ));
    InMux I__477 (
            .O(N__3039),
            .I(N__3036));
    LocalMux I__476 (
            .O(N__3036),
            .I(N__3033));
    Span12Mux_h I__475 (
            .O(N__3033),
            .I(N__3030));
    Span12Mux_v I__474 (
            .O(N__3030),
            .I(N__3027));
    Odrv12 I__473 (
            .O(N__3027),
            .I(consolereset_c));
    InMux I__472 (
            .O(N__3024),
            .I(N__3021));
    LocalMux I__471 (
            .O(N__3021),
            .I(N__3018));
    Span4Mux_h I__470 (
            .O(N__3018),
            .I(N__3015));
    Sp12to4 I__469 (
            .O(N__3015),
            .I(N__3012));
    Span12Mux_v I__468 (
            .O(N__3012),
            .I(N__3009));
    Span12Mux_v I__467 (
            .O(N__3009),
            .I(N__3006));
    Odrv12 I__466 (
            .O(N__3006),
            .I(altreset_c));
    CascadeMux I__465 (
            .O(N__3003),
            .I(\debounceconsolereset.out_RNOZ0Z_0_cascade_ ));
    InMux I__464 (
            .O(N__3000),
            .I(N__2997));
    LocalMux I__463 (
            .O(N__2997),
            .I(clock_out_RNIR6ER));
    CascadeMux I__462 (
            .O(N__2994),
            .I(clock_out_RNIR6ER_cascade_));
    InMux I__461 (
            .O(N__2991),
            .I(N__2988));
    LocalMux I__460 (
            .O(N__2988),
            .I(N__2983));
    InMux I__459 (
            .O(N__2987),
            .I(N__2978));
    InMux I__458 (
            .O(N__2986),
            .I(N__2978));
    Span4Mux_v I__457 (
            .O(N__2983),
            .I(N__2958));
    LocalMux I__456 (
            .O(N__2978),
            .I(N__2958));
    InMux I__455 (
            .O(N__2977),
            .I(N__2951));
    InMux I__454 (
            .O(N__2976),
            .I(N__2951));
    InMux I__453 (
            .O(N__2975),
            .I(N__2951));
    InMux I__452 (
            .O(N__2974),
            .I(N__2942));
    InMux I__451 (
            .O(N__2973),
            .I(N__2942));
    InMux I__450 (
            .O(N__2972),
            .I(N__2942));
    InMux I__449 (
            .O(N__2971),
            .I(N__2942));
    InMux I__448 (
            .O(N__2970),
            .I(N__2939));
    InMux I__447 (
            .O(N__2969),
            .I(N__2936));
    InMux I__446 (
            .O(N__2968),
            .I(N__2929));
    InMux I__445 (
            .O(N__2967),
            .I(N__2929));
    InMux I__444 (
            .O(N__2966),
            .I(N__2929));
    InMux I__443 (
            .O(N__2965),
            .I(N__2922));
    InMux I__442 (
            .O(N__2964),
            .I(N__2922));
    InMux I__441 (
            .O(N__2963),
            .I(N__2922));
    Span4Mux_h I__440 (
            .O(N__2958),
            .I(N__2919));
    LocalMux I__439 (
            .O(N__2951),
            .I(arses_counter8));
    LocalMux I__438 (
            .O(N__2942),
            .I(arses_counter8));
    LocalMux I__437 (
            .O(N__2939),
            .I(arses_counter8));
    LocalMux I__436 (
            .O(N__2936),
            .I(arses_counter8));
    LocalMux I__435 (
            .O(N__2929),
            .I(arses_counter8));
    LocalMux I__434 (
            .O(N__2922),
            .I(arses_counter8));
    Odrv4 I__433 (
            .O(N__2919),
            .I(arses_counter8));
    InMux I__432 (
            .O(N__2904),
            .I(N__2900));
    CascadeMux I__431 (
            .O(N__2903),
            .I(N__2896));
    LocalMux I__430 (
            .O(N__2900),
            .I(N__2890));
    InMux I__429 (
            .O(N__2899),
            .I(N__2887));
    InMux I__428 (
            .O(N__2896),
            .I(N__2884));
    InMux I__427 (
            .O(N__2895),
            .I(N__2877));
    InMux I__426 (
            .O(N__2894),
            .I(N__2877));
    InMux I__425 (
            .O(N__2893),
            .I(N__2877));
    Span4Mux_h I__424 (
            .O(N__2890),
            .I(N__2874));
    LocalMux I__423 (
            .O(N__2887),
            .I(slowclk));
    LocalMux I__422 (
            .O(N__2884),
            .I(slowclk));
    LocalMux I__421 (
            .O(N__2877),
            .I(slowclk));
    Odrv4 I__420 (
            .O(N__2874),
            .I(slowclk));
    CascadeMux I__419 (
            .O(N__2865),
            .I(N__2862));
    InMux I__418 (
            .O(N__2862),
            .I(N__2859));
    LocalMux I__417 (
            .O(N__2859),
            .I(\dig2.m54_am ));
    IoInMux I__416 (
            .O(N__2856),
            .I(N__2853));
    LocalMux I__415 (
            .O(N__2853),
            .I(N__2850));
    Span12Mux_s4_v I__414 (
            .O(N__2850),
            .I(N__2847));
    Span12Mux_v I__413 (
            .O(N__2847),
            .I(N__2844));
    Odrv12 I__412 (
            .O(N__2844),
            .I(leds_1_i_0_1));
    InMux I__411 (
            .O(N__2841),
            .I(N__2838));
    LocalMux I__410 (
            .O(N__2838),
            .I(\dig2.m75_ns_1 ));
    InMux I__409 (
            .O(N__2835),
            .I(N__2832));
    LocalMux I__408 (
            .O(N__2832),
            .I(\dig2.m69_am ));
    CascadeMux I__407 (
            .O(N__2829),
            .I(N__2826));
    InMux I__406 (
            .O(N__2826),
            .I(N__2823));
    LocalMux I__405 (
            .O(N__2823),
            .I(\dig2.m69_bm ));
    IoInMux I__404 (
            .O(N__2820),
            .I(N__2817));
    LocalMux I__403 (
            .O(N__2817),
            .I(N__2814));
    IoSpan4Mux I__402 (
            .O(N__2814),
            .I(N__2811));
    IoSpan4Mux I__401 (
            .O(N__2811),
            .I(N__2808));
    Sp12to4 I__400 (
            .O(N__2808),
            .I(N__2805));
    Span12Mux_s6_v I__399 (
            .O(N__2805),
            .I(N__2802));
    Odrv12 I__398 (
            .O(N__2802),
            .I(leds_1_i_0_2));
    InMux I__397 (
            .O(N__2799),
            .I(N__2796));
    LocalMux I__396 (
            .O(N__2796),
            .I(\dig2.N_78 ));
    CascadeMux I__395 (
            .O(N__2793),
            .I(N__2790));
    InMux I__394 (
            .O(N__2790),
            .I(N__2787));
    LocalMux I__393 (
            .O(N__2787),
            .I(\dig2.N_76 ));
    IoInMux I__392 (
            .O(N__2784),
            .I(N__2781));
    LocalMux I__391 (
            .O(N__2781),
            .I(N__2778));
    IoSpan4Mux I__390 (
            .O(N__2778),
            .I(N__2775));
    Span4Mux_s2_v I__389 (
            .O(N__2775),
            .I(N__2772));
    Span4Mux_h I__388 (
            .O(N__2772),
            .I(N__2769));
    Sp12to4 I__387 (
            .O(N__2769),
            .I(N__2766));
    Span12Mux_v I__386 (
            .O(N__2766),
            .I(N__2763));
    Odrv12 I__385 (
            .O(N__2763),
            .I(leds_1_i_0_3));
    CascadeMux I__384 (
            .O(N__2760),
            .I(\dig2.m39_ns_1_cascade_ ));
    InMux I__383 (
            .O(N__2757),
            .I(N__2754));
    LocalMux I__382 (
            .O(N__2754),
            .I(\dig2.N_40 ));
    InMux I__381 (
            .O(N__2751),
            .I(N__2748));
    LocalMux I__380 (
            .O(N__2748),
            .I(\dig2.i3_mux ));
    InMux I__379 (
            .O(N__2745),
            .I(N__2742));
    LocalMux I__378 (
            .O(N__2742),
            .I(\dig2.N_59 ));
    InMux I__377 (
            .O(N__2739),
            .I(N__2736));
    LocalMux I__376 (
            .O(N__2736),
            .I(\dig2.leds_17_i_ns_1_2 ));
    InMux I__375 (
            .O(N__2733),
            .I(N__2730));
    LocalMux I__374 (
            .O(N__2730),
            .I(\dig2.m18_am ));
    IoInMux I__373 (
            .O(N__2727),
            .I(N__2724));
    LocalMux I__372 (
            .O(N__2724),
            .I(N__2721));
    IoSpan4Mux I__371 (
            .O(N__2721),
            .I(N__2718));
    Sp12to4 I__370 (
            .O(N__2718),
            .I(N__2715));
    Span12Mux_v I__369 (
            .O(N__2715),
            .I(N__2712));
    Span12Mux_h I__368 (
            .O(N__2712),
            .I(N__2709));
    Odrv12 I__367 (
            .O(N__2709),
            .I(leds_1_i_3));
    InMux I__366 (
            .O(N__2706),
            .I(N__2703));
    LocalMux I__365 (
            .O(N__2703),
            .I(\dig2.m13_bm ));
    InMux I__364 (
            .O(N__2700),
            .I(N__2697));
    LocalMux I__363 (
            .O(N__2697),
            .I(\dig2.N_42 ));
    InMux I__362 (
            .O(N__2694),
            .I(N__2690));
    InMux I__361 (
            .O(N__2693),
            .I(N__2687));
    LocalMux I__360 (
            .O(N__2690),
            .I(\arses.counterZ0Z_11 ));
    LocalMux I__359 (
            .O(N__2687),
            .I(\arses.counterZ0Z_11 ));
    InMux I__358 (
            .O(N__2682),
            .I(N__2678));
    InMux I__357 (
            .O(N__2681),
            .I(N__2675));
    LocalMux I__356 (
            .O(N__2678),
            .I(\arses.counterZ0Z_10 ));
    LocalMux I__355 (
            .O(N__2675),
            .I(\arses.counterZ0Z_10 ));
    CascadeMux I__354 (
            .O(N__2670),
            .I(\arses.un1_counterlt11_cascade_ ));
    InMux I__353 (
            .O(N__2667),
            .I(N__2663));
    InMux I__352 (
            .O(N__2666),
            .I(N__2660));
    LocalMux I__351 (
            .O(N__2663),
            .I(\arses.counterZ0Z_9 ));
    LocalMux I__350 (
            .O(N__2660),
            .I(\arses.counterZ0Z_9 ));
    InMux I__349 (
            .O(N__2655),
            .I(N__2651));
    InMux I__348 (
            .O(N__2654),
            .I(N__2648));
    LocalMux I__347 (
            .O(N__2651),
            .I(\arses.counterZ0Z_14 ));
    LocalMux I__346 (
            .O(N__2648),
            .I(\arses.counterZ0Z_14 ));
    InMux I__345 (
            .O(N__2643),
            .I(N__2639));
    InMux I__344 (
            .O(N__2642),
            .I(N__2636));
    LocalMux I__343 (
            .O(N__2639),
            .I(\arses.counterZ0Z_13 ));
    LocalMux I__342 (
            .O(N__2636),
            .I(\arses.counterZ0Z_13 ));
    CascadeMux I__341 (
            .O(N__2631),
            .I(\arses.un1_counterlt13_0_cascade_ ));
    InMux I__340 (
            .O(N__2628),
            .I(N__2624));
    InMux I__339 (
            .O(N__2627),
            .I(N__2621));
    LocalMux I__338 (
            .O(N__2624),
            .I(\arses.counterZ0Z_12 ));
    LocalMux I__337 (
            .O(N__2621),
            .I(\arses.counterZ0Z_12 ));
    CascadeMux I__336 (
            .O(N__2616),
            .I(arses_counter8_cascade_));
    IoInMux I__335 (
            .O(N__2613),
            .I(N__2610));
    LocalMux I__334 (
            .O(N__2610),
            .I(N__2607));
    Span4Mux_s2_v I__333 (
            .O(N__2607),
            .I(N__2604));
    Span4Mux_v I__332 (
            .O(N__2604),
            .I(N__2601));
    Odrv4 I__331 (
            .O(N__2601),
            .I(\arses.clock_out_RNIR6ERZ0Z_0 ));
    CascadeMux I__330 (
            .O(N__2598),
            .I(N__2595));
    InMux I__329 (
            .O(N__2595),
            .I(N__2592));
    LocalMux I__328 (
            .O(N__2592),
            .I(N__2587));
    InMux I__327 (
            .O(N__2591),
            .I(N__2582));
    InMux I__326 (
            .O(N__2590),
            .I(N__2582));
    Odrv4 I__325 (
            .O(N__2587),
            .I(\arses.counterZ0Z_1 ));
    LocalMux I__324 (
            .O(N__2582),
            .I(\arses.counterZ0Z_1 ));
    InMux I__323 (
            .O(N__2577),
            .I(N__2571));
    InMux I__322 (
            .O(N__2576),
            .I(N__2568));
    InMux I__321 (
            .O(N__2575),
            .I(N__2563));
    InMux I__320 (
            .O(N__2574),
            .I(N__2563));
    LocalMux I__319 (
            .O(N__2571),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__318 (
            .O(N__2568),
            .I(\arses.counterZ0Z_0 ));
    LocalMux I__317 (
            .O(N__2563),
            .I(\arses.counterZ0Z_0 ));
    IoInMux I__316 (
            .O(N__2556),
            .I(N__2553));
    LocalMux I__315 (
            .O(N__2553),
            .I(N__2550));
    Odrv4 I__314 (
            .O(N__2550),
            .I(lcol3_c));
    CascadeMux I__313 (
            .O(N__2547),
            .I(\dig2.m13_am_cascade_ ));
    InMux I__312 (
            .O(N__2544),
            .I(N__2541));
    LocalMux I__311 (
            .O(N__2541),
            .I(\dig2.leds_17_i_0_ns_1_1 ));
    InMux I__310 (
            .O(N__2538),
            .I(N__2534));
    InMux I__309 (
            .O(N__2537),
            .I(N__2531));
    LocalMux I__308 (
            .O(N__2534),
            .I(\debounceup.counterZ0Z_3 ));
    LocalMux I__307 (
            .O(N__2531),
            .I(\debounceup.counterZ0Z_3 ));
    CascadeMux I__306 (
            .O(N__2526),
            .I(\debounceup.counter19_2_cascade_ ));
    InMux I__305 (
            .O(N__2523),
            .I(N__2520));
    LocalMux I__304 (
            .O(N__2520),
            .I(\debounceup.counter_RNO_0_0_2 ));
    CascadeMux I__303 (
            .O(N__2517),
            .I(\debounceup.counter19_cascade_ ));
    InMux I__302 (
            .O(N__2514),
            .I(N__2510));
    InMux I__301 (
            .O(N__2513),
            .I(N__2507));
    LocalMux I__300 (
            .O(N__2510),
            .I(\debounceup.counterZ0Z_2 ));
    LocalMux I__299 (
            .O(N__2507),
            .I(\debounceup.counterZ0Z_2 ));
    InMux I__298 (
            .O(N__2502),
            .I(N__2492));
    InMux I__297 (
            .O(N__2501),
            .I(N__2492));
    InMux I__296 (
            .O(N__2500),
            .I(N__2492));
    InMux I__295 (
            .O(N__2499),
            .I(N__2489));
    LocalMux I__294 (
            .O(N__2492),
            .I(N__2486));
    LocalMux I__293 (
            .O(N__2489),
            .I(\debounceup.counterZ0Z_4 ));
    Odrv4 I__292 (
            .O(N__2486),
            .I(\debounceup.counterZ0Z_4 ));
    InMux I__291 (
            .O(N__2481),
            .I(N__2476));
    InMux I__290 (
            .O(N__2480),
            .I(N__2471));
    InMux I__289 (
            .O(N__2479),
            .I(N__2471));
    LocalMux I__288 (
            .O(N__2476),
            .I(\debounceup.counter19_2 ));
    LocalMux I__287 (
            .O(N__2471),
            .I(\debounceup.counter19_2 ));
    CascadeMux I__286 (
            .O(N__2466),
            .I(\dig2.m18_bm_cascade_ ));
    IoInMux I__285 (
            .O(N__2463),
            .I(N__2460));
    LocalMux I__284 (
            .O(N__2460),
            .I(N__2457));
    Span4Mux_s2_v I__283 (
            .O(N__2457),
            .I(N__2454));
    Span4Mux_v I__282 (
            .O(N__2454),
            .I(N__2451));
    Span4Mux_v I__281 (
            .O(N__2451),
            .I(N__2448));
    Span4Mux_v I__280 (
            .O(N__2448),
            .I(N__2445));
    Odrv4 I__279 (
            .O(N__2445),
            .I(leds_1_i_1));
    InMux I__278 (
            .O(N__2442),
            .I(N__2438));
    InMux I__277 (
            .O(N__2441),
            .I(N__2435));
    LocalMux I__276 (
            .O(N__2438),
            .I(\arses.counterZ0Z_7 ));
    LocalMux I__275 (
            .O(N__2435),
            .I(\arses.counterZ0Z_7 ));
    InMux I__274 (
            .O(N__2430),
            .I(N__2426));
    InMux I__273 (
            .O(N__2429),
            .I(N__2423));
    LocalMux I__272 (
            .O(N__2426),
            .I(\arses.counterZ0Z_6 ));
    LocalMux I__271 (
            .O(N__2423),
            .I(\arses.counterZ0Z_6 ));
    CascadeMux I__270 (
            .O(N__2418),
            .I(N__2415));
    InMux I__269 (
            .O(N__2415),
            .I(N__2411));
    InMux I__268 (
            .O(N__2414),
            .I(N__2408));
    LocalMux I__267 (
            .O(N__2411),
            .I(N__2405));
    LocalMux I__266 (
            .O(N__2408),
            .I(\arses.counterZ0Z_5 ));
    Odrv4 I__265 (
            .O(N__2405),
            .I(\arses.counterZ0Z_5 ));
    InMux I__264 (
            .O(N__2400),
            .I(N__2396));
    InMux I__263 (
            .O(N__2399),
            .I(N__2393));
    LocalMux I__262 (
            .O(N__2396),
            .I(\arses.counterZ0Z_8 ));
    LocalMux I__261 (
            .O(N__2393),
            .I(\arses.counterZ0Z_8 ));
    InMux I__260 (
            .O(N__2388),
            .I(N__2384));
    InMux I__259 (
            .O(N__2387),
            .I(N__2381));
    LocalMux I__258 (
            .O(N__2384),
            .I(\arses.counterZ0Z_3 ));
    LocalMux I__257 (
            .O(N__2381),
            .I(\arses.counterZ0Z_3 ));
    InMux I__256 (
            .O(N__2376),
            .I(N__2372));
    InMux I__255 (
            .O(N__2375),
            .I(N__2369));
    LocalMux I__254 (
            .O(N__2372),
            .I(\arses.counterZ0Z_2 ));
    LocalMux I__253 (
            .O(N__2369),
            .I(\arses.counterZ0Z_2 ));
    InMux I__252 (
            .O(N__2364),
            .I(N__2360));
    InMux I__251 (
            .O(N__2363),
            .I(N__2357));
    LocalMux I__250 (
            .O(N__2360),
            .I(\arses.counterZ0Z_4 ));
    LocalMux I__249 (
            .O(N__2357),
            .I(\arses.counterZ0Z_4 ));
    CascadeMux I__248 (
            .O(N__2352),
            .I(\arses.un1_counterlto4_2_cascade_ ));
    InMux I__247 (
            .O(N__2349),
            .I(N__2346));
    LocalMux I__246 (
            .O(N__2346),
            .I(\arses.un1_counterlto8_2 ));
    InMux I__245 (
            .O(N__2343),
            .I(\arses.un2_counter_cry_7 ));
    InMux I__244 (
            .O(N__2340),
            .I(bfn_15_24_0_));
    InMux I__243 (
            .O(N__2337),
            .I(\arses.un2_counter_cry_9 ));
    InMux I__242 (
            .O(N__2334),
            .I(\arses.un2_counter_cry_10 ));
    InMux I__241 (
            .O(N__2331),
            .I(\arses.un2_counter_cry_11 ));
    InMux I__240 (
            .O(N__2328),
            .I(\arses.un2_counter_cry_12 ));
    InMux I__239 (
            .O(N__2325),
            .I(\arses.un2_counter_cry_13 ));
    IoInMux I__238 (
            .O(N__2322),
            .I(N__2319));
    LocalMux I__237 (
            .O(N__2319),
            .I(N__2316));
    IoSpan4Mux I__236 (
            .O(N__2316),
            .I(N__2313));
    Span4Mux_s1_v I__235 (
            .O(N__2313),
            .I(N__2310));
    Span4Mux_h I__234 (
            .O(N__2310),
            .I(N__2307));
    Odrv4 I__233 (
            .O(N__2307),
            .I(lcol4_c));
    IoInMux I__232 (
            .O(N__2304),
            .I(N__2301));
    LocalMux I__231 (
            .O(N__2301),
            .I(N__2298));
    IoSpan4Mux I__230 (
            .O(N__2298),
            .I(N__2295));
    Odrv4 I__229 (
            .O(N__2295),
            .I(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO));
    InMux I__228 (
            .O(N__2292),
            .I(\debounceup.un3_counter_1_cry_2 ));
    InMux I__227 (
            .O(N__2289),
            .I(\debounceup.un3_counter_1_cry_3 ));
    InMux I__226 (
            .O(N__2286),
            .I(\arses.un2_counter_cry_1 ));
    InMux I__225 (
            .O(N__2283),
            .I(\arses.un2_counter_cry_2 ));
    InMux I__224 (
            .O(N__2280),
            .I(\arses.un2_counter_cry_3 ));
    InMux I__223 (
            .O(N__2277),
            .I(\arses.un2_counter_cry_4 ));
    InMux I__222 (
            .O(N__2274),
            .I(\arses.un2_counter_cry_5 ));
    InMux I__221 (
            .O(N__2271),
            .I(\arses.un2_counter_cry_6 ));
    IoInMux I__220 (
            .O(N__2268),
            .I(N__2265));
    LocalMux I__219 (
            .O(N__2265),
            .I(N__2262));
    IoSpan4Mux I__218 (
            .O(N__2262),
            .I(N__2259));
    Span4Mux_s2_v I__217 (
            .O(N__2259),
            .I(N__2256));
    Sp12to4 I__216 (
            .O(N__2256),
            .I(N__2253));
    Span12Mux_s10_v I__215 (
            .O(N__2253),
            .I(N__2250));
    Span12Mux_v I__214 (
            .O(N__2250),
            .I(N__2247));
    Span12Mux_h I__213 (
            .O(N__2247),
            .I(N__2244));
    Odrv12 I__212 (
            .O(N__2244),
            .I(\arse.divseven.io_0_D_IN_0 ));
    IoInMux I__211 (
            .O(N__2241),
            .I(N__2238));
    LocalMux I__210 (
            .O(N__2238),
            .I(N__2235));
    Odrv4 I__209 (
            .O(N__2235),
            .I(masterreset_c_i));
    InMux I__208 (
            .O(N__2232),
            .I(\debounceup.un3_counter_1_cry_1 ));
    ClkMux I__207 (
            .O(N__2229),
            .I(N__2226));
    GlobalMux I__206 (
            .O(N__2226),
            .I(N__2223));
    gio2CtrlBuf I__205 (
            .O(N__2223),
            .I(\arse.un1_io_0_1_g ));
    IoInMux I__204 (
            .O(N__2220),
            .I(N__2217));
    LocalMux I__203 (
            .O(N__2217),
            .I(N__2214));
    IoSpan4Mux I__202 (
            .O(N__2214),
            .I(N__2211));
    Span4Mux_s3_h I__201 (
            .O(N__2211),
            .I(N__2208));
    Span4Mux_h I__200 (
            .O(N__2208),
            .I(N__2205));
    Sp12to4 I__199 (
            .O(N__2205),
            .I(N__2202));
    Span12Mux_h I__198 (
            .O(N__2202),
            .I(N__2199));
    Span12Mux_v I__197 (
            .O(N__2199),
            .I(N__2196));
    Odrv12 I__196 (
            .O(N__2196),
            .I(\top_pll_nrtthrth.PLLOUTCORE ));
    INV \INVarse.divseven.dout_0C  (
            .O(\INVarse.divseven.dout_0C_net ),
            .I(N__5740));
    INV \INVarse.apuresetoutregC  (
            .O(\INVarse.apuresetoutregC_net ),
            .I(N__5747));
    INV \INVarse.apusynclatchedC  (
            .O(\INVarse.apusynclatchedC_net ),
            .I(N__2229));
    INV \INVarse.diveight.dout_0C  (
            .O(\INVarse.diveight.dout_0C_net ),
            .I(N__5749));
    INV \INVarse.cpuclkresetC  (
            .O(\INVarse.cpuclkresetC_net ),
            .I(N__5745));
    INV \INVarse.cpuresetoutregC  (
            .O(\INVarse.cpuresetoutregC_net ),
            .I(N__5751));
    INV \INVarse.cpuresetcount_0C  (
            .O(\INVarse.cpuresetcount_0C_net ),
            .I(N__5750));
    defparam IN_MUX_bfv_27_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_27_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_27_10_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_24_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_17_0_));
    defparam IN_MUX_bfv_20_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_17_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\arses.un2_counter_cry_8 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_29_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_29_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_29_7_0_));
    ICE_GB \arses.clock_out_RNIR6ER_1  (
            .USERSIGNALTOGLOBALBUFFER(N__2613),
            .GLOBALBUFFEROUTPUT(N_111_g));
    ICE_GB \top_pll_nrtthrth.PLLOUTCORE_derived_clock_RNIRGL5  (
            .USERSIGNALTOGLOBALBUFFER(N__2220),
            .GLOBALBUFFEROUTPUT(PLLOUTCORE_g));
    ICE_GB \arse.divseven.io_0_RNIIG08  (
            .USERSIGNALTOGLOBALBUFFER(N__2268),
            .GLOBALBUFFEROUTPUT(\arse.un1_io_0_1_g ));
    ICE_GB masterreset_ibuf_RNIKP26_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2241),
            .GLOBALBUFFEROUTPUT(masterreset_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam masterreset_ibuf_RNIKP26_LC_3_16_6.C_ON=1'b0;
    defparam masterreset_ibuf_RNIKP26_LC_3_16_6.SEQ_MODE=4'b0000;
    defparam masterreset_ibuf_RNIKP26_LC_3_16_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 masterreset_ibuf_RNIKP26_LC_3_16_6 (
            .in0(N__4871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(masterreset_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.un3_counter_1_cry_1_c_LC_15_18_0 .C_ON=1'b1;
    defparam \debounceup.un3_counter_1_cry_1_c_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \debounceup.un3_counter_1_cry_1_c_LC_15_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debounceup.un3_counter_1_cry_1_c_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__3320),
            .in2(N__3347),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\debounceup.un3_counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_RNO_0_2_LC_15_18_1 .C_ON=1'b1;
    defparam \debounceup.counter_RNO_0_2_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \debounceup.counter_RNO_0_2_LC_15_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \debounceup.counter_RNO_0_2_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__2514),
            .in2(_gnd_net_),
            .in3(N__2232),
            .lcout(\debounceup.counter_RNO_0_0_2 ),
            .ltout(),
            .carryin(\debounceup.un3_counter_1_cry_1 ),
            .carryout(\debounceup.un3_counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_3_LC_15_18_2 .C_ON=1'b1;
    defparam \debounceup.counter_3_LC_15_18_2 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_3_LC_15_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \debounceup.counter_3_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__2538),
            .in2(_gnd_net_),
            .in3(N__2292),
            .lcout(\debounceup.counterZ0Z_3 ),
            .ltout(),
            .carryin(\debounceup.un3_counter_1_cry_2 ),
            .carryout(\debounceup.un3_counter_1_cry_3 ),
            .clk(N__4492),
            .ce(N__4596),
            .sr(_gnd_net_));
    defparam \debounceup.counter_4_LC_15_18_3 .C_ON=1'b0;
    defparam \debounceup.counter_4_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_4_LC_15_18_3 .LUT_INIT=16'b0000010100001000;
    LogicCell40 \debounceup.counter_4_LC_15_18_3  (
            .in0(N__2499),
            .in1(N__2481),
            .in2(N__4652),
            .in3(N__2289),
            .lcout(\debounceup.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4492),
            .ce(N__4596),
            .sr(_gnd_net_));
    defparam \arses.un2_counter_cry_1_c_LC_15_23_0 .C_ON=1'b1;
    defparam \arses.un2_counter_cry_1_c_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \arses.un2_counter_cry_1_c_LC_15_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \arses.un2_counter_cry_1_c_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__2576),
            .in2(N__2598),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\arses.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_2_LC_15_23_1 .C_ON=1'b1;
    defparam \arses.counter_2_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_2_LC_15_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_2_LC_15_23_1  (
            .in0(N__2971),
            .in1(N__2376),
            .in2(_gnd_net_),
            .in3(N__2286),
            .lcout(\arses.counterZ0Z_2 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_1 ),
            .carryout(\arses.un2_counter_cry_2 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_3_LC_15_23_2 .C_ON=1'b1;
    defparam \arses.counter_3_LC_15_23_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_3_LC_15_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_3_LC_15_23_2  (
            .in0(N__2963),
            .in1(N__2388),
            .in2(_gnd_net_),
            .in3(N__2283),
            .lcout(\arses.counterZ0Z_3 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_2 ),
            .carryout(\arses.un2_counter_cry_3 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_4_LC_15_23_3 .C_ON=1'b1;
    defparam \arses.counter_4_LC_15_23_3 .SEQ_MODE=4'b1001;
    defparam \arses.counter_4_LC_15_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_4_LC_15_23_3  (
            .in0(N__2972),
            .in1(N__2364),
            .in2(_gnd_net_),
            .in3(N__2280),
            .lcout(\arses.counterZ0Z_4 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_3 ),
            .carryout(\arses.un2_counter_cry_4 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_5_LC_15_23_4 .C_ON=1'b1;
    defparam \arses.counter_5_LC_15_23_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_5_LC_15_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_5_LC_15_23_4  (
            .in0(N__2964),
            .in1(N__2414),
            .in2(_gnd_net_),
            .in3(N__2277),
            .lcout(\arses.counterZ0Z_5 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_4 ),
            .carryout(\arses.un2_counter_cry_5 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_6_LC_15_23_5 .C_ON=1'b1;
    defparam \arses.counter_6_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_6_LC_15_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_6_LC_15_23_5  (
            .in0(N__2973),
            .in1(N__2430),
            .in2(_gnd_net_),
            .in3(N__2274),
            .lcout(\arses.counterZ0Z_6 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_5 ),
            .carryout(\arses.un2_counter_cry_6 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_7_LC_15_23_6 .C_ON=1'b1;
    defparam \arses.counter_7_LC_15_23_6 .SEQ_MODE=4'b1000;
    defparam \arses.counter_7_LC_15_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_7_LC_15_23_6  (
            .in0(N__2965),
            .in1(N__2442),
            .in2(_gnd_net_),
            .in3(N__2271),
            .lcout(\arses.counterZ0Z_7 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_6 ),
            .carryout(\arses.un2_counter_cry_7 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_8_LC_15_23_7 .C_ON=1'b1;
    defparam \arses.counter_8_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \arses.counter_8_LC_15_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_8_LC_15_23_7  (
            .in0(N__2974),
            .in1(N__2400),
            .in2(_gnd_net_),
            .in3(N__2343),
            .lcout(\arses.counterZ0Z_8 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_7 ),
            .carryout(\arses.un2_counter_cry_8 ),
            .clk(N__4506),
            .ce(),
            .sr(N__4048));
    defparam \arses.counter_9_LC_15_24_0 .C_ON=1'b1;
    defparam \arses.counter_9_LC_15_24_0 .SEQ_MODE=4'b1000;
    defparam \arses.counter_9_LC_15_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_9_LC_15_24_0  (
            .in0(N__2968),
            .in1(N__2667),
            .in2(_gnd_net_),
            .in3(N__2340),
            .lcout(\arses.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\arses.un2_counter_cry_9 ),
            .clk(N__4509),
            .ce(),
            .sr(N__4049));
    defparam \arses.counter_10_LC_15_24_1 .C_ON=1'b1;
    defparam \arses.counter_10_LC_15_24_1 .SEQ_MODE=4'b1000;
    defparam \arses.counter_10_LC_15_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_10_LC_15_24_1  (
            .in0(N__2975),
            .in1(N__2682),
            .in2(_gnd_net_),
            .in3(N__2337),
            .lcout(\arses.counterZ0Z_10 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_9 ),
            .carryout(\arses.un2_counter_cry_10 ),
            .clk(N__4509),
            .ce(),
            .sr(N__4049));
    defparam \arses.counter_11_LC_15_24_2 .C_ON=1'b1;
    defparam \arses.counter_11_LC_15_24_2 .SEQ_MODE=4'b1000;
    defparam \arses.counter_11_LC_15_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_11_LC_15_24_2  (
            .in0(N__2966),
            .in1(N__2694),
            .in2(_gnd_net_),
            .in3(N__2334),
            .lcout(\arses.counterZ0Z_11 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_10 ),
            .carryout(\arses.un2_counter_cry_11 ),
            .clk(N__4509),
            .ce(),
            .sr(N__4049));
    defparam \arses.counter_12_LC_15_24_3 .C_ON=1'b1;
    defparam \arses.counter_12_LC_15_24_3 .SEQ_MODE=4'b1000;
    defparam \arses.counter_12_LC_15_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_12_LC_15_24_3  (
            .in0(N__2976),
            .in1(N__2628),
            .in2(_gnd_net_),
            .in3(N__2331),
            .lcout(\arses.counterZ0Z_12 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_11 ),
            .carryout(\arses.un2_counter_cry_12 ),
            .clk(N__4509),
            .ce(),
            .sr(N__4049));
    defparam \arses.counter_13_LC_15_24_4 .C_ON=1'b1;
    defparam \arses.counter_13_LC_15_24_4 .SEQ_MODE=4'b1000;
    defparam \arses.counter_13_LC_15_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_13_LC_15_24_4  (
            .in0(N__2967),
            .in1(N__2643),
            .in2(_gnd_net_),
            .in3(N__2328),
            .lcout(\arses.counterZ0Z_13 ),
            .ltout(),
            .carryin(\arses.un2_counter_cry_12 ),
            .carryout(\arses.un2_counter_cry_13 ),
            .clk(N__4509),
            .ce(),
            .sr(N__4049));
    defparam \arses.counter_14_LC_15_24_5 .C_ON=1'b0;
    defparam \arses.counter_14_LC_15_24_5 .SEQ_MODE=4'b1000;
    defparam \arses.counter_14_LC_15_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \arses.counter_14_LC_15_24_5  (
            .in0(N__2977),
            .in1(N__2655),
            .in2(_gnd_net_),
            .in3(N__2325),
            .lcout(\arses.counterZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4509),
            .ce(),
            .sr(N__4049));
    defparam lcolreg_3_LC_15_31_0.C_ON=1'b0;
    defparam lcolreg_3_LC_15_31_0.SEQ_MODE=4'b1000;
    defparam lcolreg_3_LC_15_31_0.LUT_INIT=16'b0101010111111111;
    LogicCell40 lcolreg_3_LC_15_31_0 (
            .in0(N__3581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3732),
            .lcout(lcol4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4512),
            .ce(N__4592),
            .sr(_gnd_net_));
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_6.C_ON=1'b0;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_PACKAGEPIN_0_c_g_THRU_LUT4_0_LC_16_1_6 (
            .in0(N__4518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_PACKAGEPIN_0_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_RNI5J0P_2_LC_16_18_0 .C_ON=1'b0;
    defparam \debounceup.counter_RNI5J0P_2_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \debounceup.counter_RNI5J0P_2_LC_16_18_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \debounceup.counter_RNI5J0P_2_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__2537),
            .in2(_gnd_net_),
            .in3(N__2513),
            .lcout(\debounceup.counter19_2 ),
            .ltout(\debounceup.counter19_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_RNIADHU1_1_LC_16_18_1 .C_ON=1'b0;
    defparam \debounceup.counter_RNIADHU1_1_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \debounceup.counter_RNIADHU1_1_LC_16_18_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \debounceup.counter_RNIADHU1_1_LC_16_18_1  (
            .in0(N__2500),
            .in1(N__3321),
            .in2(N__2526),
            .in3(N__3342),
            .lcout(\debounceup.counter19 ),
            .ltout(\debounceup.counter19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_2_LC_16_18_2 .C_ON=1'b0;
    defparam \debounceup.counter_2_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_2_LC_16_18_2 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \debounceup.counter_2_LC_16_18_2  (
            .in0(N__2480),
            .in1(N__2523),
            .in2(N__2517),
            .in3(N__2502),
            .lcout(\debounceup.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4489),
            .ce(N__4595),
            .sr(_gnd_net_));
    defparam \debounceup.counter_0_LC_16_18_3 .C_ON=1'b0;
    defparam \debounceup.counter_0_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_0_LC_16_18_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \debounceup.counter_0_LC_16_18_3  (
            .in0(N__2501),
            .in1(N__2479),
            .in2(_gnd_net_),
            .in3(N__3343),
            .lcout(\debounceup.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4489),
            .ce(N__4595),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m18_bm_LC_16_18_6 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m18_bm_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m18_bm_LC_16_18_6 .LUT_INIT=16'b1101010110001010;
    LogicCell40 \dig2.leds_cnst_3_1__m18_bm_LC_16_18_6  (
            .in0(N__4414),
            .in1(N__3572),
            .in2(N__4321),
            .in3(N__3095),
            .lcout(),
            .ltout(\dig2.m18_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_1_LC_16_18_7 .C_ON=1'b0;
    defparam \dig2.leds_1_i_1_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_1_LC_16_18_7 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \dig2.leds_1_i_1_LC_16_18_7  (
            .in0(N__4190),
            .in1(N__2733),
            .in2(N__2466),
            .in3(N__2544),
            .lcout(leds_1_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4489),
            .ce(N__4595),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIA58_5_LC_16_23_1 .C_ON=1'b0;
    defparam \arses.counter_RNIA58_5_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIA58_5_LC_16_23_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \arses.counter_RNIA58_5_LC_16_23_1  (
            .in0(N__2441),
            .in1(N__2429),
            .in2(N__2418),
            .in3(N__2399),
            .lcout(\arses.un1_counterlto8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI1L5_2_LC_16_23_2 .C_ON=1'b0;
    defparam \arses.counter_RNI1L5_2_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI1L5_2_LC_16_23_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \arses.counter_RNI1L5_2_LC_16_23_2  (
            .in0(N__2387),
            .in1(N__2375),
            .in2(_gnd_net_),
            .in3(N__2574),
            .lcout(),
            .ltout(\arses.un1_counterlto4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOKH_1_LC_16_23_3 .C_ON=1'b0;
    defparam \arses.counter_RNIOKH_1_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOKH_1_LC_16_23_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \arses.counter_RNIOKH_1_LC_16_23_3  (
            .in0(N__2363),
            .in1(N__2590),
            .in2(N__2352),
            .in3(N__2349),
            .lcout(),
            .ltout(\arses.un1_counterlt11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNI04C4_9_LC_16_23_4 .C_ON=1'b0;
    defparam \arses.counter_RNI04C4_9_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNI04C4_9_LC_16_23_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \arses.counter_RNI04C4_9_LC_16_23_4  (
            .in0(N__2693),
            .in1(N__2681),
            .in2(N__2670),
            .in3(N__2666),
            .lcout(),
            .ltout(\arses.un1_counterlt13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_RNIOS0A_14_LC_16_23_5 .C_ON=1'b0;
    defparam \arses.counter_RNIOS0A_14_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \arses.counter_RNIOS0A_14_LC_16_23_5 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \arses.counter_RNIOS0A_14_LC_16_23_5  (
            .in0(N__2654),
            .in1(N__2642),
            .in2(N__2631),
            .in3(N__2627),
            .lcout(arses_counter8),
            .ltout(arses_counter8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_0_LC_16_23_6 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_0_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_0_LC_16_23_6 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \arses.clock_out_RNIR6ER_0_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(N__4834),
            .in2(N__2616),
            .in3(N__2904),
            .lcout(\arses.clock_out_RNIR6ERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.counter_1_LC_16_23_7 .C_ON=1'b0;
    defparam \arses.counter_1_LC_16_23_7 .SEQ_MODE=4'b1001;
    defparam \arses.counter_1_LC_16_23_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \arses.counter_1_LC_16_23_7  (
            .in0(N__2575),
            .in1(N__2970),
            .in2(_gnd_net_),
            .in3(N__2591),
            .lcout(\arses.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4503),
            .ce(),
            .sr(N__4050));
    defparam \arses.counter_0_LC_16_24_7 .C_ON=1'b0;
    defparam \arses.counter_0_LC_16_24_7 .SEQ_MODE=4'b1001;
    defparam \arses.counter_0_LC_16_24_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \arses.counter_0_LC_16_24_7  (
            .in0(_gnd_net_),
            .in1(N__2969),
            .in2(_gnd_net_),
            .in3(N__2577),
            .lcout(\arses.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4507),
            .ce(),
            .sr(N__4052));
    defparam lcolreg_2_LC_16_31_3.C_ON=1'b0;
    defparam lcolreg_2_LC_16_31_3.SEQ_MODE=4'b1000;
    defparam lcolreg_2_LC_16_31_3.LUT_INIT=16'b1111111100110011;
    LogicCell40 lcolreg_2_LC_16_31_3 (
            .in0(_gnd_net_),
            .in1(N__3739),
            .in2(_gnd_net_),
            .in3(N__3571),
            .lcout(lcol3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4511),
            .ce(N__4591),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m13_am_LC_17_18_1 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m13_am_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m13_am_LC_17_18_1 .LUT_INIT=16'b1000101001111010;
    LogicCell40 \dig2.leds_cnst_3_1__m13_am_LC_17_18_1  (
            .in0(N__4412),
            .in1(N__3721),
            .in2(N__4311),
            .in3(N__3552),
            .lcout(),
            .ltout(\dig2.m13_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_1_LC_17_18_2 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_1_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_1_LC_17_18_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_1_LC_17_18_2  (
            .in0(N__4181),
            .in1(N__4119),
            .in2(N__2547),
            .in3(N__2706),
            .lcout(\dig2.leds_17_i_0_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m18_am_LC_17_18_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m18_am_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m18_am_LC_17_18_4 .LUT_INIT=16'b0000001000000100;
    LogicCell40 \dig2.leds_cnst_3_1__m18_am_LC_17_18_4  (
            .in0(N__3553),
            .in1(N__4299),
            .in2(N__3738),
            .in3(N__4413),
            .lcout(\dig2.m18_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m77_LC_18_16_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m77_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m77_LC_18_16_7 .LUT_INIT=16'b0101101100111111;
    LogicCell40 \dig2.leds_cnst_3_1__m77_LC_18_16_7  (
            .in0(N__5615),
            .in1(N__3725),
            .in2(N__5315),
            .in3(N__3554),
            .lcout(\dig2.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_3_LC_18_17_3 .C_ON=1'b0;
    defparam \dig2.leds_1_i_3_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_3_LC_18_17_3 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \dig2.leds_1_i_3_LC_18_17_3  (
            .in0(N__2700),
            .in1(N__4194),
            .in2(N__4110),
            .in3(N__2757),
            .lcout(leds_1_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4487),
            .ce(N__4597),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m61_LC_18_18_2 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m61_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m61_LC_18_18_2 .LUT_INIT=16'b0101101110100000;
    LogicCell40 \dig2.leds_cnst_3_1__m61_LC_18_18_2  (
            .in0(N__5609),
            .in1(N__3659),
            .in2(N__5312),
            .in3(N__3476),
            .lcout(\dig2.i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m58_LC_18_18_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m58_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m58_LC_18_18_4 .LUT_INIT=16'b0000001110000100;
    LogicCell40 \dig2.leds_cnst_3_1__m58_LC_18_18_4  (
            .in0(N__5610),
            .in1(N__3660),
            .in2(N__5311),
            .in3(N__3477),
            .lcout(\dig2.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m13_bm_LC_18_18_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m13_bm_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m13_bm_LC_18_18_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \dig2.leds_cnst_3_1__m13_bm_LC_18_18_7  (
            .in0(N__3478),
            .in1(N__4403),
            .in2(N__4295),
            .in3(N__3666),
            .lcout(\dig2.m13_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m41_LC_19_16_1 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m41_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m41_LC_19_16_1 .LUT_INIT=16'b0101100101111111;
    LogicCell40 \dig2.leds_cnst_3_1__m41_LC_19_16_1  (
            .in0(N__4384),
            .in1(N__3559),
            .in2(N__4322),
            .in3(N__3687),
            .lcout(\dig2.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m75_ns_LC_19_16_2 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m75_ns_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m75_ns_LC_19_16_2 .LUT_INIT=16'b0011000001010101;
    LogicCell40 \dig2.leds_cnst_3_1__m75_ns_LC_19_16_2  (
            .in0(N__2841),
            .in1(N__4996),
            .in2(N__3096),
            .in3(N__5614),
            .lcout(\dig2.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m54_am_LC_19_16_5 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m54_am_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m54_am_LC_19_16_5 .LUT_INIT=16'b0000000001000010;
    LogicCell40 \dig2.leds_cnst_3_1__m54_am_LC_19_16_5  (
            .in0(N__5611),
            .in1(N__3558),
            .in2(N__5313),
            .in3(N__3686),
            .lcout(\dig2.m54_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m69_am_LC_19_16_6 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m69_am_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m69_am_LC_19_16_6 .LUT_INIT=16'b1100101001100111;
    LogicCell40 \dig2.leds_cnst_3_1__m69_am_LC_19_16_6  (
            .in0(N__3560),
            .in1(N__5613),
            .in2(N__3720),
            .in3(N__5293),
            .lcout(\dig2.m69_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m69_bm_LC_19_16_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m69_bm_LC_19_16_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m69_bm_LC_19_16_7 .LUT_INIT=16'b1001001111000100;
    LogicCell40 \dig2.leds_cnst_3_1__m69_bm_LC_19_16_7  (
            .in0(N__5612),
            .in1(N__3561),
            .in2(N__5314),
            .in3(N__3691),
            .lcout(\dig2.m69_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_2_LC_19_17_1 .C_ON=1'b0;
    defparam \dig1.leds_1_i_2_LC_19_17_1 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_2_LC_19_17_1 .LUT_INIT=16'b1101100001010101;
    LogicCell40 \dig1.leds_1_i_2_LC_19_17_1  (
            .in0(N__2739),
            .in1(N__2835),
            .in2(N__2829),
            .in3(N__5689),
            .lcout(leds_1_i_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4490),
            .ce(N__4598),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_0_LC_19_17_4 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_0_LC_19_17_4 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_0_LC_19_17_4 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \debounceconsolereset.counter_0_LC_19_17_4  (
            .in0(N__3196),
            .in1(N__3182),
            .in2(_gnd_net_),
            .in3(N__3137),
            .lcout(\debounceconsolereset.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4490),
            .ce(N__4598),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_1_LC_19_17_5 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_1_LC_19_17_5 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_1_LC_19_17_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \debounceconsolereset.counter_1_LC_19_17_5  (
            .in0(N__3138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3161),
            .lcout(\debounceconsolereset.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4490),
            .ce(N__4598),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_2_LC_19_17_6 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_2_LC_19_17_6 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_2_LC_19_17_6 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \debounceconsolereset.counter_2_LC_19_17_6  (
            .in0(N__3240),
            .in1(N__3183),
            .in2(N__3201),
            .in3(N__3113),
            .lcout(\debounceconsolereset.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4490),
            .ce(N__4598),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_3_LC_19_17_7 .C_ON=1'b0;
    defparam \dig1.leds_1_i_3_LC_19_17_7 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_3_LC_19_17_7 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \dig1.leds_1_i_3_LC_19_17_7  (
            .in0(N__2799),
            .in1(N__5690),
            .in2(N__2793),
            .in3(N__4997),
            .lcout(leds_1_i_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4490),
            .ce(N__4598),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m39_ns_1_LC_19_18_3 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m39_ns_1_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m39_ns_1_LC_19_18_3 .LUT_INIT=16'b0111010111110101;
    LogicCell40 \dig2.leds_cnst_3_1__m39_ns_1_LC_19_18_3  (
            .in0(N__4375),
            .in1(N__3658),
            .in2(N__4118),
            .in3(N__3475),
            .lcout(),
            .ltout(\dig2.m39_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m39_ns_LC_19_18_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m39_ns_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m39_ns_LC_19_18_4 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \dig2.leds_cnst_3_1__m39_ns_LC_19_18_4  (
            .in0(N__4323),
            .in1(N__4114),
            .in2(N__2760),
            .in3(N__3087),
            .lcout(\dig2.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_18_5 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_18_5 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \dig2.leds_cnst_3_1__leds_17_i_ns_1_2_LC_19_18_5  (
            .in0(N__2751),
            .in1(N__4995),
            .in2(N__5691),
            .in3(N__2745),
            .lcout(\dig2.leds_17_i_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m3_LC_19_18_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m3_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m3_LC_19_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dig2.leds_cnst_3_1__m3_LC_19_18_7  (
            .in0(_gnd_net_),
            .in1(N__3657),
            .in2(_gnd_net_),
            .in3(N__3474),
            .lcout(col_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam col_1_LC_19_19_0.C_ON=1'b0;
    defparam col_1_LC_19_19_0.SEQ_MODE=4'b1000;
    defparam col_1_LC_19_19_0.LUT_INIT=16'b1100110010101100;
    LogicCell40 col_1_LC_19_19_0 (
            .in0(N__3091),
            .in1(N__3672),
            .in2(N__2903),
            .in3(N__3000),
            .lcout(colZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4495),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_RNO_0_LC_19_19_3 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNO_0_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNO_0_LC_19_19_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \debounceconsolereset.out_RNO_0_LC_19_19_3  (
            .in0(N__2894),
            .in1(N__3112),
            .in2(N__4864),
            .in3(N__2987),
            .lcout(),
            .ltout(\debounceconsolereset.out_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.out_LC_19_19_4 .C_ON=1'b0;
    defparam \debounceconsolereset.out_LC_19_19_4 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.out_LC_19_19_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \debounceconsolereset.out_LC_19_19_4  (
            .in0(N__3039),
            .in1(N__3024),
            .in2(N__3003),
            .in3(N__5387),
            .lcout(debouncedconsolereset),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4495),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_RNIR6ER_LC_19_19_6 .C_ON=1'b0;
    defparam \arses.clock_out_RNIR6ER_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \arses.clock_out_RNIR6ER_LC_19_19_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \arses.clock_out_RNIR6ER_LC_19_19_6  (
            .in0(N__2986),
            .in1(N__4853),
            .in2(_gnd_net_),
            .in3(N__2893),
            .lcout(clock_out_RNIR6ER),
            .ltout(clock_out_RNIR6ER_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam col_0_LC_19_19_7.C_ON=1'b0;
    defparam col_0_LC_19_19_7.SEQ_MODE=4'b1000;
    defparam col_0_LC_19_19_7.LUT_INIT=16'b1111010100001010;
    LogicCell40 col_0_LC_19_19_7 (
            .in0(N__2895),
            .in1(_gnd_net_),
            .in2(N__2994),
            .in3(N__3508),
            .lcout(colZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4495),
            .ce(),
            .sr(_gnd_net_));
    defparam \arses.clock_out_LC_19_20_2 .C_ON=1'b0;
    defparam \arses.clock_out_LC_19_20_2 .SEQ_MODE=4'b1000;
    defparam \arses.clock_out_LC_19_20_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \arses.clock_out_LC_19_20_2  (
            .in0(N__2991),
            .in1(N__4863),
            .in2(_gnd_net_),
            .in3(N__2899),
            .lcout(slowclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4500),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig1.leds_1_i_1_LC_20_16_3 .C_ON=1'b0;
    defparam \dig1.leds_1_i_1_LC_20_16_3 .SEQ_MODE=4'b1000;
    defparam \dig1.leds_1_i_1_LC_20_16_3 .LUT_INIT=16'b1011001110010001;
    LogicCell40 \dig1.leds_1_i_1_LC_20_16_3  (
            .in0(N__5688),
            .in1(N__3048),
            .in2(N__2865),
            .in3(N__3057),
            .lcout(leds_1_i_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4491),
            .ce(N__4601),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m75_ns_1_LC_20_16_6 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m75_ns_1_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m75_ns_1_LC_20_16_6 .LUT_INIT=16'b0111010111110101;
    LogicCell40 \dig2.leds_cnst_3_1__m75_ns_1_LC_20_16_6  (
            .in0(N__5283),
            .in1(N__3692),
            .in2(N__4994),
            .in3(N__3557),
            .lcout(\dig2.m75_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.un3_counter_1_cry_1_c_LC_20_17_0 .C_ON=1'b1;
    defparam \debounceconsolereset.un3_counter_1_cry_1_c_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.un3_counter_1_cry_1_c_LC_20_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debounceconsolereset.un3_counter_1_cry_1_c_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(N__3136),
            .in2(N__3162),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_17_0_),
            .carryout(\debounceconsolereset.un3_counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNO_0_2_LC_20_17_1 .C_ON=1'b1;
    defparam \debounceconsolereset.counter_RNO_0_2_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNO_0_2_LC_20_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \debounceconsolereset.counter_RNO_0_2_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(N__3213),
            .in2(_gnd_net_),
            .in3(N__3234),
            .lcout(\debounceconsolereset.counter_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_1_cry_1 ),
            .carryout(\debounceconsolereset.un3_counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_3_LC_20_17_2 .C_ON=1'b1;
    defparam \debounceconsolereset.counter_3_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_3_LC_20_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \debounceconsolereset.counter_3_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(N__3225),
            .in2(_gnd_net_),
            .in3(N__3231),
            .lcout(\debounceconsolereset.counterZ0Z_3 ),
            .ltout(),
            .carryin(\debounceconsolereset.un3_counter_1_cry_2 ),
            .carryout(\debounceconsolereset.un3_counter_1_cry_3 ),
            .clk(N__4493),
            .ce(N__4600),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_4_LC_20_17_3 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_4_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \debounceconsolereset.counter_4_LC_20_17_3 .LUT_INIT=16'b0000001100001000;
    LogicCell40 \debounceconsolereset.counter_4_LC_20_17_3  (
            .in0(N__3200),
            .in1(N__3181),
            .in2(N__3117),
            .in3(N__3228),
            .lcout(\debounceconsolereset.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4493),
            .ce(N__4600),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNI7OV8_2_LC_20_18_0 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_RNI7OV8_2_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNI7OV8_2_LC_20_18_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \debounceconsolereset.counter_RNI7OV8_2_LC_20_18_0  (
            .in0(_gnd_net_),
            .in1(N__3224),
            .in2(_gnd_net_),
            .in3(N__3212),
            .lcout(\debounceconsolereset.counter19_2 ),
            .ltout(\debounceconsolereset.counter19_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceconsolereset.counter_RNIV9FM_1_LC_20_18_1 .C_ON=1'b0;
    defparam \debounceconsolereset.counter_RNIV9FM_1_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.counter_RNIV9FM_1_LC_20_18_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \debounceconsolereset.counter_RNIV9FM_1_LC_20_18_1  (
            .in0(N__3180),
            .in1(N__3157),
            .in2(N__3141),
            .in3(N__3135),
            .lcout(\debounceconsolereset.counter19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m54_bm_LC_20_18_2 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m54_bm_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m54_bm_LC_20_18_2 .LUT_INIT=16'b1000111111010000;
    LogicCell40 \dig2.leds_cnst_3_1__m54_bm_LC_20_18_2  (
            .in0(N__5616),
            .in1(N__3488),
            .in2(N__5325),
            .in3(N__3086),
            .lcout(\dig2.m54_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_0_LC_21_14_6.C_ON=1'b0;
    defparam delayConstant_0_LC_21_14_6.SEQ_MODE=4'b1000;
    defparam delayConstant_0_LC_21_14_6.LUT_INIT=16'b0101010110011001;
    LogicCell40 delayConstant_0_LC_21_14_6 (
            .in0(N__5282),
            .in1(N__4719),
            .in2(_gnd_net_),
            .in3(N__4758),
            .lcout(delayConstantZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4488),
            .ce(),
            .sr(N__4051));
    defparam \dig2.leds_cnst_3_1__leds_17_i_ns_1_1_LC_21_16_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__leds_17_i_ns_1_1_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__leds_17_i_ns_1_1_LC_21_16_4 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \dig2.leds_cnst_3_1__leds_17_i_ns_1_1_LC_21_16_4  (
            .in0(N__4998),
            .in1(N__3294),
            .in2(N__5683),
            .in3(N__3288),
            .lcout(\dig2.leds_17_i_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.counter_1_LC_21_19_0 .C_ON=1'b0;
    defparam \debounceup.counter_1_LC_21_19_0 .SEQ_MODE=4'b1000;
    defparam \debounceup.counter_1_LC_21_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounceup.counter_1_LC_21_19_0  (
            .in0(_gnd_net_),
            .in1(N__3351),
            .in2(_gnd_net_),
            .in3(N__3313),
            .lcout(\debounceup.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4501),
            .ce(N__4599),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m49_bm_LC_22_15_2 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m49_bm_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m49_bm_LC_22_15_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \dig2.leds_cnst_3_1__m49_bm_LC_22_15_2  (
            .in0(N__5586),
            .in1(N__3709),
            .in2(N__3586),
            .in3(N__5239),
            .lcout(\dig2.m49_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m33_am_LC_22_15_3 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m33_am_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m33_am_LC_22_15_3 .LUT_INIT=16'b1101001010011011;
    LogicCell40 \dig2.leds_cnst_3_1__m33_am_LC_22_15_3  (
            .in0(N__3579),
            .in1(N__4415),
            .in2(N__4303),
            .in3(N__3719),
            .lcout(\dig2.m33_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m49_am_LC_22_15_6 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m49_am_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m49_am_LC_22_15_6 .LUT_INIT=16'b1101011100001010;
    LogicCell40 \dig2.leds_cnst_3_1__m49_am_LC_22_15_6  (
            .in0(N__5587),
            .in1(N__3710),
            .in2(N__3587),
            .in3(N__5238),
            .lcout(\dig2.m49_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m33_bm_LC_22_16_0 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m33_bm_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m33_bm_LC_22_16_0 .LUT_INIT=16'b1010010000111100;
    LogicCell40 \dig2.leds_cnst_3_1__m33_bm_LC_22_16_0  (
            .in0(N__4416),
            .in1(N__3737),
            .in2(N__3580),
            .in3(N__4294),
            .lcout(),
            .ltout(\dig2.m33_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_1_i_2_LC_22_16_1 .C_ON=1'b0;
    defparam \dig2.leds_1_i_2_LC_22_16_1 .SEQ_MODE=4'b1000;
    defparam \dig2.leds_1_i_2_LC_22_16_1 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \dig2.leds_1_i_2_LC_22_16_1  (
            .in0(N__4185),
            .in1(N__3282),
            .in2(N__3276),
            .in3(N__3252),
            .lcout(leds_1_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4496),
            .ce(N__4603),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m22_LC_23_17_4 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m22_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m22_LC_23_17_4 .LUT_INIT=16'b0001000110000100;
    LogicCell40 \dig2.leds_cnst_3_1__m22_LC_23_17_4  (
            .in0(N__4404),
            .in1(N__3736),
            .in2(N__4304),
            .in3(N__3556),
            .lcout(),
            .ltout(\dig2.N_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_23_17_5 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_23_17_5 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \dig2.leds_cnst_3_1__leds_17_i_0_ns_1_2_LC_23_17_5  (
            .in0(N__3246),
            .in1(N__4186),
            .in2(N__3255),
            .in3(N__4109),
            .lcout(\dig2.leds_17_i_0_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dig2.leds_cnst_3_1__m25_LC_23_17_7 .C_ON=1'b0;
    defparam \dig2.leds_cnst_3_1__m25_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \dig2.leds_cnst_3_1__m25_LC_23_17_7 .LUT_INIT=16'b0110011010001010;
    LogicCell40 \dig2.leds_cnst_3_1__m25_LC_23_17_7  (
            .in0(N__3555),
            .in1(N__4405),
            .in2(N__3745),
            .in3(N__4285),
            .lcout(\dig2.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_0_LC_23_18_2 .C_ON=1'b0;
    defparam \debouncedn.counter_0_LC_23_18_2 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_0_LC_23_18_2 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \debouncedn.counter_0_LC_23_18_2  (
            .in0(N__3980),
            .in1(N__3956),
            .in2(_gnd_net_),
            .in3(N__3930),
            .lcout(\debouncedn.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4504),
            .ce(N__4602),
            .sr(_gnd_net_));
    defparam lcolreg_0_LC_23_30_3.C_ON=1'b0;
    defparam lcolreg_0_LC_23_30_3.SEQ_MODE=4'b1000;
    defparam lcolreg_0_LC_23_30_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 lcolreg_0_LC_23_30_3 (
            .in0(_gnd_net_),
            .in1(N__3752),
            .in2(_gnd_net_),
            .in3(N__3591),
            .lcout(lcol1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4513),
            .ce(N__4594),
            .sr(_gnd_net_));
    defparam lcolreg_1_LC_23_31_7.C_ON=1'b0;
    defparam lcolreg_1_LC_23_31_7.SEQ_MODE=4'b1000;
    defparam lcolreg_1_LC_23_31_7.LUT_INIT=16'b1100110011111111;
    LogicCell40 lcolreg_1_LC_23_31_7 (
            .in0(_gnd_net_),
            .in1(N__3753),
            .in2(_gnd_net_),
            .in3(N__3582),
            .lcout(lcol2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4514),
            .ce(N__4593),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_RNIVDIV_2_LC_24_16_2 .C_ON=1'b0;
    defparam \debouncedn.counter_RNIVDIV_2_LC_24_16_2 .SEQ_MODE=4'b0000;
    defparam \debouncedn.counter_RNIVDIV_2_LC_24_16_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \debouncedn.counter_RNIVDIV_2_LC_24_16_2  (
            .in0(_gnd_net_),
            .in1(N__3365),
            .in2(_gnd_net_),
            .in3(N__3386),
            .lcout(\debouncedn.counter19_2 ),
            .ltout(\debouncedn.counter19_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_RNIB0UE2_1_LC_24_16_3 .C_ON=1'b0;
    defparam \debouncedn.counter_RNIB0UE2_1_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \debouncedn.counter_RNIB0UE2_1_LC_24_16_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \debouncedn.counter_RNIB0UE2_1_LC_24_16_3  (
            .in0(N__3954),
            .in1(N__3933),
            .in2(N__3393),
            .in3(N__3903),
            .lcout(\debouncedn.counter19 ),
            .ltout(\debouncedn.counter19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_2_LC_24_16_4 .C_ON=1'b0;
    defparam \debouncedn.counter_2_LC_24_16_4 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_2_LC_24_16_4 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \debouncedn.counter_2_LC_24_16_4  (
            .in0(N__3957),
            .in1(N__3375),
            .in2(N__3390),
            .in3(N__3979),
            .lcout(\debouncedn.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4502),
            .ce(N__4606),
            .sr(_gnd_net_));
    defparam \debouncedn.un3_counter_1_cry_1_c_LC_24_17_0 .C_ON=1'b1;
    defparam \debouncedn.un3_counter_1_cry_1_c_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \debouncedn.un3_counter_1_cry_1_c_LC_24_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \debouncedn.un3_counter_1_cry_1_c_LC_24_17_0  (
            .in0(_gnd_net_),
            .in1(N__3898),
            .in2(N__3932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_24_17_0_),
            .carryout(\debouncedn.un3_counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_RNO_0_2_LC_24_17_1 .C_ON=1'b1;
    defparam \debouncedn.counter_RNO_0_2_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \debouncedn.counter_RNO_0_2_LC_24_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \debouncedn.counter_RNO_0_2_LC_24_17_1  (
            .in0(_gnd_net_),
            .in1(N__3387),
            .in2(_gnd_net_),
            .in3(N__3369),
            .lcout(\debouncedn.counter_RNO_0_1_2 ),
            .ltout(),
            .carryin(\debouncedn.un3_counter_1_cry_1 ),
            .carryout(\debouncedn.un3_counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_3_LC_24_17_2 .C_ON=1'b1;
    defparam \debouncedn.counter_3_LC_24_17_2 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_3_LC_24_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \debouncedn.counter_3_LC_24_17_2  (
            .in0(_gnd_net_),
            .in1(N__3366),
            .in2(_gnd_net_),
            .in3(N__3354),
            .lcout(\debouncedn.counterZ0Z_3 ),
            .ltout(),
            .carryin(\debouncedn.un3_counter_1_cry_2 ),
            .carryout(\debouncedn.un3_counter_1_cry_3 ),
            .clk(N__4505),
            .ce(N__4605),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_4_LC_24_17_3 .C_ON=1'b0;
    defparam \debouncedn.counter_4_LC_24_17_3 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_4_LC_24_17_3 .LUT_INIT=16'b0001000100100000;
    LogicCell40 \debouncedn.counter_4_LC_24_17_3  (
            .in0(N__3955),
            .in1(N__3878),
            .in2(N__3984),
            .in3(N__3960),
            .lcout(\debouncedn.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4505),
            .ce(N__4605),
            .sr(_gnd_net_));
    defparam \debouncedn.counter_1_LC_24_18_4 .C_ON=1'b0;
    defparam \debouncedn.counter_1_LC_24_18_4 .SEQ_MODE=4'b1000;
    defparam \debouncedn.counter_1_LC_24_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debouncedn.counter_1_LC_24_18_4  (
            .in0(_gnd_net_),
            .in1(N__3931),
            .in2(_gnd_net_),
            .in3(N__3902),
            .lcout(\debouncedn.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4508),
            .ce(N__4604),
            .sr(_gnd_net_));
    defparam \debouncedn.out_LC_26_12_6 .C_ON=1'b0;
    defparam \debouncedn.out_LC_26_12_6 .SEQ_MODE=4'b1000;
    defparam \debouncedn.out_LC_26_12_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \debouncedn.out_LC_26_12_6  (
            .in0(N__3882),
            .in1(N__3864),
            .in2(N__4023),
            .in3(N__4614),
            .lcout(debounceddn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4497),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_26_25_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_26_25_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_26_25_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_26_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_0_c_LC_27_10_0.C_ON=1'b1;
    defparam un1_delayConstant_cry_0_c_LC_27_10_0.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_0_c_LC_27_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_delayConstant_cry_0_c_LC_27_10_0 (
            .in0(_gnd_net_),
            .in1(N__4776),
            .in2(N__5326),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_27_10_0_),
            .carryout(un1_delayConstant_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delayConstant_1_LC_27_10_1.C_ON=1'b1;
    defparam delayConstant_1_LC_27_10_1.SEQ_MODE=4'b1000;
    defparam delayConstant_1_LC_27_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_1_LC_27_10_1 (
            .in0(_gnd_net_),
            .in1(N__4002),
            .in2(N__5571),
            .in3(N__3777),
            .lcout(delayConstantZ0Z_1),
            .ltout(),
            .carryin(un1_delayConstant_cry_0),
            .carryout(un1_delayConstant_cry_1),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam delayConstant_2_LC_27_10_2.C_ON=1'b1;
    defparam delayConstant_2_LC_27_10_2.SEQ_MODE=4'b1000;
    defparam delayConstant_2_LC_27_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_2_LC_27_10_2 (
            .in0(_gnd_net_),
            .in1(N__4764),
            .in2(N__5649),
            .in3(N__3774),
            .lcout(delayConstantZ0Z_2),
            .ltout(),
            .carryin(un1_delayConstant_cry_1),
            .carryout(un1_delayConstant_cry_2),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam delayConstant_3_LC_27_10_3.C_ON=1'b1;
    defparam delayConstant_3_LC_27_10_3.SEQ_MODE=4'b1000;
    defparam delayConstant_3_LC_27_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_3_LC_27_10_3 (
            .in0(_gnd_net_),
            .in1(N__4665),
            .in2(N__4971),
            .in3(N__3771),
            .lcout(delayConstantZ0Z_3),
            .ltout(),
            .carryin(un1_delayConstant_cry_2),
            .carryout(un1_delayConstant_cry_3),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam delayConstant_4_LC_27_10_4.C_ON=1'b1;
    defparam delayConstant_4_LC_27_10_4.SEQ_MODE=4'b1000;
    defparam delayConstant_4_LC_27_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_4_LC_27_10_4 (
            .in0(_gnd_net_),
            .in1(N__3996),
            .in2(N__4374),
            .in3(N__4326),
            .lcout(delayConstantZ0Z_4),
            .ltout(),
            .carryin(un1_delayConstant_cry_3),
            .carryout(un1_delayConstant_cry_4),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam delayConstant_5_LC_27_10_5.C_ON=1'b1;
    defparam delayConstant_5_LC_27_10_5.SEQ_MODE=4'b1000;
    defparam delayConstant_5_LC_27_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_5_LC_27_10_5 (
            .in0(_gnd_net_),
            .in1(N__3990),
            .in2(N__4259),
            .in3(N__4197),
            .lcout(delayConstantZ0Z_5),
            .ltout(),
            .carryin(un1_delayConstant_cry_4),
            .carryout(un1_delayConstant_cry_5),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam delayConstant_6_LC_27_10_6.C_ON=1'b1;
    defparam delayConstant_6_LC_27_10_6.SEQ_MODE=4'b1000;
    defparam delayConstant_6_LC_27_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delayConstant_6_LC_27_10_6 (
            .in0(_gnd_net_),
            .in1(N__4770),
            .in2(N__4171),
            .in3(N__4125),
            .lcout(delayConstantZ0Z_6),
            .ltout(),
            .carryin(un1_delayConstant_cry_5),
            .carryout(un1_delayConstant_cry_6),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam delayConstant_7_LC_27_10_7.C_ON=1'b0;
    defparam delayConstant_7_LC_27_10_7.SEQ_MODE=4'b1000;
    defparam delayConstant_7_LC_27_10_7.LUT_INIT=16'b1000011101111000;
    LogicCell40 delayConstant_7_LC_27_10_7 (
            .in0(N__4706),
            .in1(N__4751),
            .in2(N__4089),
            .in3(N__4122),
            .lcout(delayConstantZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4494),
            .ce(),
            .sr(N__4053));
    defparam olddn_LC_27_11_0.C_ON=1'b0;
    defparam olddn_LC_27_11_0.SEQ_MODE=4'b1000;
    defparam olddn_LC_27_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 olddn_LC_27_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4019),
            .lcout(olddnZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4498),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIEENH_LC_27_11_2.C_ON=1'b0;
    defparam olddn_RNIEENH_LC_27_11_2.SEQ_MODE=4'b0000;
    defparam olddn_RNIEENH_LC_27_11_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 olddn_RNIEENH_LC_27_11_2 (
            .in0(_gnd_net_),
            .in1(N__4029),
            .in2(_gnd_net_),
            .in3(N__4018),
            .lcout(olddn_RNIEENHZ0),
            .ltout(olddn_RNIEENHZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_0_LC_27_11_3.C_ON=1'b0;
    defparam olddn_RNIM5BH1_0_LC_27_11_3.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_0_LC_27_11_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 olddn_RNIM5BH1_0_LC_27_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4005),
            .in3(N__4694),
            .lcout(olddn_RNIM5BH1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_3_LC_28_10_0.C_ON=1'b0;
    defparam olddn_RNIM5BH1_3_LC_28_10_0.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_3_LC_28_10_0.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNIM5BH1_3_LC_28_10_0 (
            .in0(N__4748),
            .in1(_gnd_net_),
            .in2(N__4711),
            .in3(_gnd_net_),
            .lcout(olddn_RNIM5BH1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_1_LC_28_10_1.C_ON=1'b0;
    defparam olddn_RNIM5BH1_1_LC_28_10_1.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_1_LC_28_10_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_1_LC_28_10_1 (
            .in0(_gnd_net_),
            .in1(N__4702),
            .in2(_gnd_net_),
            .in3(N__4749),
            .lcout(olddn_RNIM5BH1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam oldup_RNI8NJV_LC_28_10_2.C_ON=1'b0;
    defparam oldup_RNI8NJV_LC_28_10_2.SEQ_MODE=4'b0000;
    defparam oldup_RNI8NJV_LC_28_10_2.LUT_INIT=16'b1111111101110111;
    LogicCell40 oldup_RNI8NJV_LC_28_10_2 (
            .in0(N__4852),
            .in1(N__4659),
            .in2(_gnd_net_),
            .in3(N__4541),
            .lcout(delayConstant17_i),
            .ltout(delayConstant17_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_delayConstant_cry_0_c_RNO_LC_28_10_3.C_ON=1'b0;
    defparam un1_delayConstant_cry_0_c_RNO_LC_28_10_3.SEQ_MODE=4'b0000;
    defparam un1_delayConstant_cry_0_c_RNO_LC_28_10_3.LUT_INIT=16'b1111111100001111;
    LogicCell40 un1_delayConstant_cry_0_c_RNO_LC_28_10_3 (
            .in0(N__5327),
            .in1(_gnd_net_),
            .in2(N__4779),
            .in3(N__4745),
            .lcout(un1_delayConstant_cry_0_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_4_LC_28_10_4.C_ON=1'b0;
    defparam olddn_RNIM5BH1_4_LC_28_10_4.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_4_LC_28_10_4.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNIM5BH1_4_LC_28_10_4 (
            .in0(N__4750),
            .in1(_gnd_net_),
            .in2(N__4712),
            .in3(_gnd_net_),
            .lcout(olddn_RNIM5BH1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_LC_28_10_5.C_ON=1'b0;
    defparam olddn_RNIM5BH1_LC_28_10_5.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_LC_28_10_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 olddn_RNIM5BH1_LC_28_10_5 (
            .in0(_gnd_net_),
            .in1(N__4695),
            .in2(_gnd_net_),
            .in3(N__4746),
            .lcout(olddn_RNIM5BHZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam olddn_RNIM5BH1_2_LC_28_10_6.C_ON=1'b0;
    defparam olddn_RNIM5BH1_2_LC_28_10_6.SEQ_MODE=4'b0000;
    defparam olddn_RNIM5BH1_2_LC_28_10_6.LUT_INIT=16'b1010000010100000;
    LogicCell40 olddn_RNIM5BH1_2_LC_28_10_6 (
            .in0(N__4747),
            .in1(_gnd_net_),
            .in2(N__4710),
            .in3(_gnd_net_),
            .lcout(olddn_RNIM5BH1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam oldup_LC_28_10_7.C_ON=1'b0;
    defparam oldup_LC_28_10_7.SEQ_MODE=4'b1000;
    defparam oldup_LC_28_10_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 oldup_LC_28_10_7 (
            .in0(N__4542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(oldupZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4499),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounceup.out_LC_28_18_5 .C_ON=1'b0;
    defparam \debounceup.out_LC_28_18_5 .SEQ_MODE=4'b1000;
    defparam \debounceup.out_LC_28_18_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \debounceup.out_LC_28_18_5  (
            .in0(N__4653),
            .in1(N__4632),
            .in2(N__4540),
            .in3(N__4613),
            .lcout(debouncedup),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4510),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_0_LC_29_7_0 .C_ON=1'b1;
    defparam \arse.cpuresetcount_0_LC_29_7_0 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_0_LC_29_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_0_LC_29_7_0  (
            .in0(_gnd_net_),
            .in1(N__5172),
            .in2(N__5481),
            .in3(N__5480),
            .lcout(\arse.cpuresetcountZ0Z_0 ),
            .ltout(),
            .carryin(bfn_29_7_0_),
            .carryout(\arse.un1_cpuresetcount_1_cry_0 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_1_LC_29_7_1 .C_ON=1'b1;
    defparam \arse.cpuresetcount_1_LC_29_7_1 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_1_LC_29_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_1_LC_29_7_1  (
            .in0(_gnd_net_),
            .in1(N__5138),
            .in2(_gnd_net_),
            .in3(N__4419),
            .lcout(\arse.cpuresetcountZ0Z_1 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_0 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_1 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_2_LC_29_7_2 .C_ON=1'b1;
    defparam \arse.cpuresetcount_2_LC_29_7_2 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_2_LC_29_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_2_LC_29_7_2  (
            .in0(_gnd_net_),
            .in1(N__5121),
            .in2(_gnd_net_),
            .in3(N__4914),
            .lcout(\arse.cpuresetcountZ0Z_2 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_1 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_2 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_3_LC_29_7_3 .C_ON=1'b1;
    defparam \arse.cpuresetcount_3_LC_29_7_3 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_3_LC_29_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_3_LC_29_7_3  (
            .in0(_gnd_net_),
            .in1(N__5055),
            .in2(_gnd_net_),
            .in3(N__4911),
            .lcout(\arse.cpuresetcountZ0Z_3 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_2 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_3 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_4_LC_29_7_4 .C_ON=1'b1;
    defparam \arse.cpuresetcount_4_LC_29_7_4 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_4_LC_29_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_4_LC_29_7_4  (
            .in0(_gnd_net_),
            .in1(N__5103),
            .in2(_gnd_net_),
            .in3(N__4908),
            .lcout(\arse.cpuresetcountZ0Z_4 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_3 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_4 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_5_LC_29_7_5 .C_ON=1'b1;
    defparam \arse.cpuresetcount_5_LC_29_7_5 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_5_LC_29_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_5_LC_29_7_5  (
            .in0(_gnd_net_),
            .in1(N__5156),
            .in2(_gnd_net_),
            .in3(N__4905),
            .lcout(\arse.cpuresetcountZ0Z_5 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_4 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_5 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_6_LC_29_7_6 .C_ON=1'b1;
    defparam \arse.cpuresetcount_6_LC_29_7_6 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_6_LC_29_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \arse.cpuresetcount_6_LC_29_7_6  (
            .in0(_gnd_net_),
            .in1(N__5067),
            .in2(_gnd_net_),
            .in3(N__4902),
            .lcout(\arse.cpuresetcountZ0Z_6 ),
            .ltout(),
            .carryin(\arse.un1_cpuresetcount_1_cry_5 ),
            .carryout(\arse.un1_cpuresetcount_1_cry_6 ),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \arse.cpuresetcount_7_LC_29_7_7 .C_ON=1'b0;
    defparam \arse.cpuresetcount_7_LC_29_7_7 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetcount_7_LC_29_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \arse.cpuresetcount_7_LC_29_7_7  (
            .in0(_gnd_net_),
            .in1(N__5079),
            .in2(_gnd_net_),
            .in3(N__4899),
            .lcout(\arse.cpuresetcountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuresetcount_0C_net ),
            .ce(),
            .sr(N__5028));
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_2 .C_ON=1'b0;
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_2 .SEQ_MODE=4'b0000;
    defparam \debounceconsolereset.out_RNI1B6C_LC_29_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \debounceconsolereset.out_RNI1B6C_LC_29_8_2  (
            .in0(N__5413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debouncedconsolereset_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_LC_30_6_2 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_LC_30_6_2 .SEQ_MODE=4'b1000;
    defparam \arse.cpuresetoutreg_LC_30_6_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \arse.cpuresetoutreg_LC_30_6_2  (
            .in0(_gnd_net_),
            .in1(N__4892),
            .in2(_gnd_net_),
            .in3(N__5085),
            .lcout(\arse.cpuresetoutregZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuresetoutregC_net ),
            .ce(),
            .sr(N__5027));
    defparam \arse.cpuclkreset_RNO_1_LC_30_7_1 .C_ON=1'b0;
    defparam \arse.cpuclkreset_RNO_1_LC_30_7_1 .SEQ_MODE=4'b0000;
    defparam \arse.cpuclkreset_RNO_1_LC_30_7_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \arse.cpuclkreset_RNO_1_LC_30_7_1  (
            .in0(N__5119),
            .in1(N__5170),
            .in2(N__5157),
            .in3(N__5134),
            .lcout(),
            .ltout(\arse.m8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuclkreset_RNO_0_LC_30_7_2 .C_ON=1'b0;
    defparam \arse.cpuclkreset_RNO_0_LC_30_7_2 .SEQ_MODE=4'b0000;
    defparam \arse.cpuclkreset_RNO_0_LC_30_7_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \arse.cpuclkreset_RNO_0_LC_30_7_2  (
            .in0(N__5469),
            .in1(N__5101),
            .in2(N__5175),
            .in3(N__5042),
            .lcout(\arse.cpuclkreset_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_1_LC_30_7_4 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_1_LC_30_7_4 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_1_LC_30_7_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \arse.cpuresetoutreg_RNO_1_LC_30_7_4  (
            .in0(N__5171),
            .in1(N__5155),
            .in2(N__5139),
            .in3(N__5120),
            .lcout(),
            .ltout(\arse.m12_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetoutreg_RNO_0_LC_30_7_5 .C_ON=1'b0;
    defparam \arse.cpuresetoutreg_RNO_0_LC_30_7_5 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetoutreg_RNO_0_LC_30_7_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \arse.cpuresetoutreg_RNO_0_LC_30_7_5  (
            .in0(N__5043),
            .in1(N__5470),
            .in2(N__5106),
            .in3(N__5102),
            .lcout(\arse.cpuresetoutreg_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuresetcount_RNIFLN61_7_LC_30_7_6 .C_ON=1'b0;
    defparam \arse.cpuresetcount_RNIFLN61_7_LC_30_7_6 .SEQ_MODE=4'b0000;
    defparam \arse.cpuresetcount_RNIFLN61_7_LC_30_7_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \arse.cpuresetcount_RNIFLN61_7_LC_30_7_6  (
            .in0(N__5078),
            .in1(N__5066),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\arse.m4_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.cpuclkreset_LC_30_8_4 .C_ON=1'b0;
    defparam \arse.cpuclkreset_LC_30_8_4 .SEQ_MODE=4'b1000;
    defparam \arse.cpuclkreset_LC_30_8_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \arse.cpuclkreset_LC_30_8_4  (
            .in0(_gnd_net_),
            .in1(N__5034),
            .in2(_gnd_net_),
            .in3(N__5516),
            .lcout(arse_cpuclkreset),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.cpuclkresetC_net ),
            .ce(),
            .sr(N__5026));
    defparam \arse.diveight.dout_0_LC_31_6_3 .C_ON=1'b0;
    defparam \arse.diveight.dout_0_LC_31_6_3 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_0_LC_31_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.diveight.dout_0_LC_31_6_3  (
            .in0(_gnd_net_),
            .in1(N__5206),
            .in2(_gnd_net_),
            .in3(N__5520),
            .lcout(\arse.diveight.doutZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.diveight.dout_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_RNI7BAS_1_LC_31_7_1 .C_ON=1'b0;
    defparam \arse.diveight.counter_RNI7BAS_1_LC_31_7_1 .SEQ_MODE=4'b0000;
    defparam \arse.diveight.counter_RNI7BAS_1_LC_31_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \arse.diveight.counter_RNI7BAS_1_LC_31_7_1  (
            .in0(_gnd_net_),
            .in1(N__5368),
            .in2(_gnd_net_),
            .in3(N__5352),
            .lcout(),
            .ltout(arse_diveight_N_123_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_2_LC_31_7_2 .C_ON=1'b0;
    defparam \arse.diveight.counter_2_LC_31_7_2 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_2_LC_31_7_2 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \arse.diveight.counter_2_LC_31_7_2  (
            .in0(N__4990),
            .in1(N__5207),
            .in2(N__4917),
            .in3(N__5514),
            .lcout(arse_diveight_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5746),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_1_LC_31_7_5 .C_ON=1'b0;
    defparam \arse.diveight.counter_1_LC_31_7_5 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_1_LC_31_7_5 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \arse.diveight.counter_1_LC_31_7_5  (
            .in0(N__5513),
            .in1(N__5369),
            .in2(N__5684),
            .in3(N__5353),
            .lcout(arse_diveight_counter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5746),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_RNO_1_LC_31_7_6 .C_ON=1'b0;
    defparam \arse.diveight.dout_RNO_1_LC_31_7_6 .SEQ_MODE=4'b0000;
    defparam \arse.diveight.dout_RNO_1_LC_31_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.diveight.dout_RNO_1_LC_31_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5512),
            .lcout(\arse.diveight.cpuclkreset_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.counter_0_LC_31_8_6 .C_ON=1'b0;
    defparam \arse.diveight.counter_0_LC_31_8_6 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.counter_0_LC_31_8_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \arse.diveight.counter_0_LC_31_8_6  (
            .in0(N__5588),
            .in1(N__5355),
            .in2(_gnd_net_),
            .in3(N__5515),
            .lcout(arse_diveight_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5742),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.apusynclatched_LC_32_3_3 .C_ON=1'b0;
    defparam \arse.apusynclatched_LC_32_3_3 .SEQ_MODE=4'b1000;
    defparam \arse.apusynclatched_LC_32_3_3 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \arse.apusynclatched_LC_32_3_3  (
            .in0(N__5487),
            .in1(N__5453),
            .in2(_gnd_net_),
            .in3(N__5424),
            .lcout(\arse.apusynclatchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.apusynclatchedC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.io_0_RNO_0_LC_32_5_0 .C_ON=1'b0;
    defparam \arse.diveight.io_0_RNO_0_LC_32_5_0 .SEQ_MODE=4'b0000;
    defparam \arse.diveight.io_0_RNO_0_LC_32_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.diveight.io_0_RNO_0_LC_32_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5442),
            .lcout(\arse.diveight.dout_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.io_0_RNO_LC_32_6_0 .C_ON=1'b0;
    defparam \arse.diveight.io_0_RNO_LC_32_6_0 .SEQ_MODE=4'b0000;
    defparam \arse.diveight.io_0_RNO_LC_32_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.diveight.io_0_RNO_LC_32_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5190),
            .lcout(\arse.diveight.dout_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.apuresetoutreg_LC_32_6_5 .C_ON=1'b0;
    defparam \arse.apuresetoutreg_LC_32_6_5 .SEQ_MODE=4'b1000;
    defparam \arse.apuresetoutreg_LC_32_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.apuresetoutreg_LC_32_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5420),
            .lcout(\arse.apuresetoutregZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.apuresetoutregC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.diveight.dout_1_LC_32_7_0 .C_ON=1'b0;
    defparam \arse.diveight.dout_1_LC_32_7_0 .SEQ_MODE=4'b1000;
    defparam \arse.diveight.dout_1_LC_32_7_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \arse.diveight.dout_1_LC_32_7_0  (
            .in0(N__5370),
            .in1(N__5354),
            .in2(N__5334),
            .in3(N__5208),
            .lcout(\arse.diveight.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5743),
            .ce(),
            .sr(N__5184));
    defparam \arse.divseven.counter_2_LC_32_8_0 .C_ON=1'b0;
    defparam \arse.divseven.counter_2_LC_32_8_0 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_2_LC_32_8_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \arse.divseven.counter_2_LC_32_8_0  (
            .in0(N__5811),
            .in1(N__5799),
            .in2(_gnd_net_),
            .in3(N__5768),
            .lcout(\arse.divseven.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5741),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_1_LC_32_8_2 .C_ON=1'b0;
    defparam \arse.divseven.counter_1_LC_32_8_2 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_1_LC_32_8_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \arse.divseven.counter_1_LC_32_8_2  (
            .in0(_gnd_net_),
            .in1(N__5810),
            .in2(_gnd_net_),
            .in3(N__5798),
            .lcout(\arse.divseven.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5741),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.counter_0_LC_32_8_4 .C_ON=1'b0;
    defparam \arse.divseven.counter_0_LC_32_8_4 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.counter_0_LC_32_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.divseven.counter_0_LC_32_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5797),
            .lcout(\arse.divseven.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5741),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_0_LC_32_9_1 .C_ON=1'b0;
    defparam \arse.divseven.dout_0_LC_32_9_1 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_0_LC_32_9_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \arse.divseven.dout_0_LC_32_9_1  (
            .in0(_gnd_net_),
            .in1(N__5767),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\arse.divseven.doutZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVarse.divseven.dout_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.io_0_RNO_0_LC_32_10_0 .C_ON=1'b0;
    defparam \arse.divseven.io_0_RNO_0_LC_32_10_0 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.io_0_RNO_0_LC_32_10_0 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \arse.divseven.io_0_RNO_0_LC_32_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5787),
            .in3(_gnd_net_),
            .lcout(\arse.divseven.dout_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.dout_1_LC_32_10_5 .C_ON=1'b0;
    defparam \arse.divseven.dout_1_LC_32_10_5 .SEQ_MODE=4'b1000;
    defparam \arse.divseven.dout_1_LC_32_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \arse.divseven.dout_1_LC_32_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5772),
            .lcout(\arse.divseven.doutZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5739),
            .ce(),
            .sr(_gnd_net_));
    defparam \arse.divseven.io_0_RNO_LC_32_10_7 .C_ON=1'b0;
    defparam \arse.divseven.io_0_RNO_LC_32_10_7 .SEQ_MODE=4'b0000;
    defparam \arse.divseven.io_0_RNO_LC_32_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \arse.divseven.io_0_RNO_LC_32_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5703),
            .lcout(\arse.divseven.dout_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
